* Spice Netlist (renamed)

*--- Top Level ---
.subckt Thermal_Camera 
.ends Thermal_Camera

