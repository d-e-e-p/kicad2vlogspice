//--- Top Level ---
module buffering_test();



endmodule

//--- Cell Definitions ---
