//--- Top Level ---
module Thermal_Camera();



endmodule

//--- Cell Definitions ---
