//--- Top Level ---
module \kicad-pyspice-example ();



endmodule

//--- Cell Definitions ---
