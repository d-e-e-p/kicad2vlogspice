* Spice Netlist (renamed)

*--- Top Level ---
.subckt ATMEGA328_Motor_Board 
.ends ATMEGA328_Motor_Board

