//--- Top Level ---
module TOP();

  wire VAL;
  wire LED0;
  wire LED1;
  wire LED2;
  wire LED3;
  wire in0;
  wire in1;
  wire in2;
  wire LED4;
  wire in3;
  wire in4;
  wire in5;
  wire LED5;

  SUB inst_sub0 (.p1(VAL), .p2(LED0));
  SUB inst_sub1 (.p1(VAL), .p2(LED0));
  SUB inst_sub2 (.p1(VAL), .p2(LED0));
  SUB inst_sub3 (.p1(VAL), .p2(LED0));
  SUB inst_sub4_0_ (.p1(VAL), .p2(LED1));
  SUB inst_sub4_1_ (.p1(VAL), .p2(LED1));
  SUB inst_sub4_2_ (.p1(VAL), .p2(LED1));
  SUB inst_sub4_3_ (.p1(VAL), .p2(LED1));
  SUB inst_sub5_0_ (.p1(VAL), .p2(LED2));
  SUB inst_sub5_1_ (.p1(VAL), .p2(LED2));
  SUB inst_sub5_2_ (.p1(VAL), .p2(LED2));
  SUB inst_sub5_3_ (.p1(VAL), .p2(LED2));
  AND U0_0_ (.p1(LED3), .p2(in0), .p3(in1), .p4(in2));
  AND U0_1_ (.p1(LED3), .p2(in0), .p3(in1), .p4(in2));
  AND U0_2_ (.p1(LED3), .p2(in0), .p3(in1), .p4(in2));
  AND U0_3_ (.p1(LED3), .p2(in0), .p3(in1), .p4(in2));
  AND unnamed_inst_0 (.p1(LED4), .p2(in3), .p3(in4), .p4(in5));
  AND unnamed_inst_1 (.p1(LED5), .p2(in3), .p3(in4), .p4(in5));

endmodule

//--- Cell Definitions ---
module TOP();
  // Stub for TOP
endmodule

module SUB();
  // Stub for SUB
endmodule

