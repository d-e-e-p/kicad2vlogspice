* Spice Netlist (renamed)

*--- Top Level ---
.subckt buffering_test 
.ends buffering_test

