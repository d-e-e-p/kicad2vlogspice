//--- Top Level ---
module \anavi-macro-pad-10 ();



endmodule

//--- Cell Definitions ---
