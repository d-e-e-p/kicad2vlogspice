* Spice Netlist (renamed)

*--- Top Level ---
.subckt kicad9_test 
.ends kicad9_test

