* Spice Netlist (renamed)

*--- Top Level ---
.subckt HDMI2USB 
.ends HDMI2USB

