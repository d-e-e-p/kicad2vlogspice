* Spice Netlist (renamed)

*--- Top Level ---
.subckt A64-OlinuXino_Rev_H 
.ends A64-OlinuXino_Rev_H

