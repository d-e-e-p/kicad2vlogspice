* Spice Netlist (renamed)

*--- Top Level ---
.subckt anavi-macro-pad-10 
.ends anavi-macro-pad-10

