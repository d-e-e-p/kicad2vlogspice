//--- Top Level ---
module components();



endmodule

//--- Cell Definitions ---
