//--- Top Level ---
module kicad9_test();



endmodule

//--- Cell Definitions ---
