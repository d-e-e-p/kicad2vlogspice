* Spice Netlist (renamed)

*--- Top Level ---
.subckt \edu-ciaa-nxp CPU_ADC0_1 CPU_ADC0_2 CPU_ADC0_3 CPU_CAN_RD CPU_CAN_TD CPU_CHJ3 CPU_DAC CPU_EECLK CPU_EECS CPU_EEDATA CPU_ENET_CRS_DV CPU_ENET_MDC CPU_ENET_MDIO CPU_ENET_REF_CLK CPU_ENET_RXD0 CPU_ENET_RXD1 CPU_ENET_TXD0 CPU_ENET_TXD1 CPU_ENET_TX_EN CPU_FT_OE CPU_FT_RST CPU_FT_TCK CPU_FT_TDI CPU_FT_TDO CPU_FT_TMS CPU_FT_TRST CPU_FT_XTIN CPU_FT_XTOUT CPU_GPIO0 CPU_GPIO1 CPU_GPIO2 CPU_GPIO3 CPU_GPIO4 CPU_GPIO5 CPU_GPIO6 CPU_GPIO7 CPU_GPIO8 CPU_I2C_SCL CPU_I2C_SDA CPU_ISP CPU_LCD1 CPU_LCD2 CPU_LCD3 CPU_LCD4 CPU_LCD_RS CPU_LED0_B CPU_LED0_G CPU_LED0_R CPU_LED1 CPU_LED2 CPU_LED3 CPU_PULS_0 CPU_PULS_1 CPU_PULS_2 CPU_PULS_3 CPU_RESET CPU_RS232_RXD CPU_RS232_TXD CPU_RS485_DIR CPU_RS485_RXD CPU_RS485_TXD CPU_RST CPU_RTCX1 CPU_RTCX2 CPU_SPI_MISO CPU_SPI_MOSI CPU_SPI_SCK CPU_TCK CPU_TDI CPU_TDO CPU_TEC_COL0 CPU_TEC_COL1 CPU_TEC_COL2 CPU_TEC_F0 CPU_TEC_F1 CPU_TEC_F2 CPU_TEC_F3 CPU_TMS CPU_TRST CPU_U2_RXD CPU_U2_TXD CPU_USB_DEBUG_VBUS CPU_USB_DM CPU_USB_DP CPU_USB_ID CPU_USB_JTAG_DM CPU_USB_JTAG_DP CPU_USB_PPWR CPU_USB_PWR_FAULT CPU_USB_VBUS CPU_XTAL1 CPU_XTAL2 CPU_nTRST GND GNDA GPIO_LCD_EN GPIO_WAKEUP USB_OTG_CHJ2 _5V _CPU_USB_JTAG_1.8V __3.3V __3.3VADC unnamed
  XH1 unnamed CONN_1
  XH2 unnamed CONN_1
  XH3 unnamed CONN_1
  XH4 unnamed CONN_1
  XF1 unnamed CONN_1
  XF2 unnamed CONN_1
  XF3 unnamed CONN_1
  XF4 unnamed CONN_1
  XF5 unnamed CONN_1
  XF6 unnamed CONN_1
  XTP1 GND CONN_1
  XU1 CPU_RS485_RXD unnamed CPU_RS485_DIR CPU_RS485_TXD GND unnamed unnamed _5V MAX3072
  XC2 _5V GND C_MINI
  XR4 _5V unnamed R_MINI
  XR7 unnamed unnamed R_MINI
  XR5 unnamed GND R_MINI
  XD1 GND unnamed ESD
  XD2 unnamed unnamed ESD
  XD3 unnamed GND ESD
  XR6 _5V unnamed R_MINI
  XR8 unnamed GND R_MINI
  XJP4 unnamed unnamed JUMPER_2
  XJP3 unnamed unnamed JUMPER_2
  XJP2 unnamed unnamed JUMPER_2
  XJ1 unnamed unnamed unnamed TB_1X3
  XR3 CPU_RS485_DIR GND R_MINI
  XR2 unnamed GND R_MINI
  XJP1 CPU_RS485_DIR unnamed JUMPER_2
  XC1 GND _5V CP_MINI
  XPS2 unnamed unnamed R
  XPS1 unnamed unnamed R
  XR9 GND unnamed R_MINI
  XR1 __3.3V CPU_RS485_RXD R_MINI
  XU2 USB_OTG_CHJ2 CPU_USB_DM CPU_USB_DP CPU_USB_VBUS PRTR5V0U2X
  XC3 CPU_USB_VBUS GND CAPAPOL
  XC4 CPU_USB_VBUS GND C
  XJ2 unnamed unnamed unnamed CPU_USB_ID GND USB_OTG_CHJ2 USB_OTG_CHJ2 USB_OTG_CHJ2 USB_OTG_CHJ2 CONN_9
  XFB2 GND USB_OTG_CHJ2 FILTER
  XFB1 unnamed CPU_USB_VBUS FILTER
  XTR1 unnamed CPU_USB_DP CPU_USB_DM unnamed TRASF_UNIP
  XU9 CPU_USB_PPWR CPU_USB_PWR_FAULT GND unnamed unnamed CPU_USB_VBUS _5V CPU_USB_VBUS MIC2025
  XC50 _5V GND C
  XR16 CPU_USB_PWR_FAULT __3.3V R
  XR17 GND CPU_USB_PPWR R
  XTH1 unnamed __3.3V THERMISTOR
  XTH2 unnamed _5V THERMISTOR
  XP1 unnamed GNDA unnamed GNDA unnamed GNDA unnamed GNDA __3.3VADC GNDA CPU_I2C_SDA unnamed GND CPU_I2C_SCL GND CPU_RS232_RXD GND CPU_RS232_TXD GND CPU_CAN_RD GND CPU_CAN_TD CPU_RESET GND CPU_TEC_COL1 GND CPU_TEC_F0 CPU_TEC_COL2 CPU_TEC_F3 CPU_TEC_F1 CPU_TEC_F2 GND CPU_TEC_COL0 GND GND CPU_ISP GPIO_WAKEUP GNDA GNDA unnamed CONN_20X2
  XP2 unnamed CPU_ENET_CRS_DV GND CPU_ENET_MDIO GND CPU_ENET_TXD0 CPU_ENET_REF_CLK CPU_ENET_TXD1 GND CPU_SPI_MISO GND unnamed CPU_SPI_SCK CPU_SPI_MOSI CPU_LCD4 GPIO_LCD_EN CPU_LCD_RS GND CPU_LCD3 GND CPU_LCD2 CPU_GPIO0 GND CPU_LCD1 CPU_GPIO2 CPU_GPIO1 CPU_GPIO4 CPU_GPIO3 CPU_GPIO6 CPU_GPIO5 GND CPU_GPIO7 GND CPU_ENET_RXD1 CPU_GPIO8 GND CPU_ENET_TX_EN GND CPU_ENET_MDC CPU_ENET_RXD0 CONN_20X2
  XR20 CPU_DAC unnamed R
  XR21 CPU_ADC0_1 unnamed R
  XR22 CPU_ADC0_2 unnamed R
  XR23 CPU_ADC0_3 unnamed R
  XTH3 unnamed __3.3V THERMISTOR
  XTH4 unnamed _5V THERMISTOR
  XC5 _5V GND CAPAPOL
  XC6 __3.3V GND CAPAPOL
  XD6 unnamed GND LED
  XR57 _5V unnamed R
  XFB3 __3.3V __3.3VADC FILTER
  XFB4 GND GNDA FILTER
  XD5 CPU_USB_DEBUG_VBUS _5V DIODESCH
  XD4 CPU_USB_VBUS _5V DIODESCH
  XU3 GND __3.3V _5V __3.3V NCP1117ST15T3G
  XC49 _5V GND C
  XZA1 GND _5V ZENER
  XD10 unnamed _5V DIODESCH
  XP4 GND unnamed CONN_2
  XC22 GND __3.3V C
  XC23 GND __3.3V C
  XC24 GND __3.3V C
  XC25 GND __3.3V C
  XC26 GND __3.3V C
  XC27 GND __3.3V C
  XC28 GND __3.3V C
  XC29 GND __3.3V C
  XC30 GND __3.3V C
  XC31 GND __3.3V C
  XC21 GND __3.3V C
  XC20 GND __3.3V C
  XC19 __3.3VADC GNDA C
  XC18 __3.3VADC GNDA C
  XR92 unnamed GND R
  XC32 __3.3VADC GNDA C
  XC33 GNDA __3.3VADC C
  XC17 unnamed GND C
  XR90 unnamed __3.3V R
  XSW5 unnamed unnamed GND GND SW_PUSH
  XR91 CPU_XTAL1 CPU_XTAL2 R
  XC14 GND CPU_XTAL1 C
  XC13 GND CPU_XTAL2 C
  XC12 GND CPU_RTCX2 C
  XC11 GND CPU_RTCX1 C
  XR98 CPU_USB_DM GND R
  XR93 unnamed __3.3V R
  XR96 CPU_USB_DP GND R
  XU4 CPU_TEC_F0 CPU_LCD2 CPU_GPIO6 CPU_GPIO7 unnamed CPU_GPIO8 CPU_LED1 CPU_LED2 CPU_LED3 __3.3V unnamed GND CPU_LCD3 unnamed __3.3V unnamed CPU_U2_TXD CPU_CAN_RD CPU_U2_RXD CPU_CAN_TD unnamed unnamed unnamed CPU_XTAL1 CPU_SPI_SCK unnamed unnamed unnamed unnamed CPU_RTCX1 CPU_RTCX2 unnamed unnamed unnamed CPU_XTAL2 GPIO_WAKEUP __3.3V CPU_TEC_COL1 CPU_TEC_COL2 CPU_ISP GNDA unnamed __3.3VADC unnamed CPU_ADC0_3 unnamed CPU_ENET_MDC __3.3V unnamed CPU_ADC0_2 unnamed CPU_LCD_RS unnamed unnamed CPU_USB_DP unnamed CPU_ADC0_1 CPU_USB_DM CPU_USB_VBUS CPU_USB_ID unnamed unnamed __3.3V CPU_TDI CPU_TCK unnamed CPU_nTRST CPU_TEC_F1 CPU_TMS CPU_TDO CPU_ENET_RXD1 GPIO_LCD_EN CPU_ENET_TX_EN CPU_LCD4 __3.3V unnamed CPU_PULS_0 unnamed GND GND __3.3V CPU_PULS_1 CPU_PULS_2 CPU_SPI_MISO unnamed unnamed CPU_SPI_MOSI CPU_TEC_COL0 CPU_PULS_3 __3.3V unnamed unnamed unnamed unnamed unnamed unnamed unnamed unnamed unnamed __3.3V CPU_DAC unnamed unnamed CPU_ENET_RXD0 unnamed CPU_ENET_CRS_DV unnamed CPU_ENET_MDIO CPU_ENET_TXD0 CPU_ENET_REF_CLK CPU_RS485_TXD CPU_TEC_F3 CPU_ENET_TXD1 __3.3V CPU_RS485_RXD unnamed CPU_GPIO0 CPU_LED0_R GND __3.3V CPU_RS485_DIR CPU_USB_PPWR CPU_TEC_F2 CPU_GPIO1 CPU_LED0_G CPU_GPIO2 CPU_USB_PWR_FAULT CPU_LED0_B CPU_GPIO3 CPU_GPIO4 CPU_RS232_TXD CPU_RS232_RXD unnamed CPU_LCD1 unnamed unnamed CPU_I2C_SCL CPU_I2C_SDA __3.3V unnamed unnamed CPU_GPIO5 unnamed unnamed LPC4337JBD144
  XP3 __3.3V CPU_RESET CPU_TMS GND CPU_TCK GND CPU_TDO unnamed CPU_TDI GND CONN_5X2
  XC16 GND CPU_FT_XTOUT C
  XC15 GND CPU_FT_XTIN C
  XU5 CPU_EECS CPU_EECLK CPU_EEDATA unnamed GND __3.3V GND __3.3V _93C56
  XC34 __3.3V GND C
  XR101 CPU_EEDATA unnamed R
  XR102 __3.3V CPU_EECS R
  XR100 __3.3V CPU_EECLK R
  XR99 __3.3V unnamed R
  XR94 CPU_nTRST __3.3V R
  XR95 __3.3V CPU_I2C_SCL R
  XR97 __3.3V CPU_I2C_SDA R
  XC48 GND __3.3V C
  XC40 GND __3.3V C
  XR105 unnamed CPU_FT_OE R
  XR106 unnamed GND R
  XR108 GND unnamed R
  XR107 GND unnamed R
  XU7 CPU_FT_TCK unnamed GND unnamed unnamed CPU_RST CPU_TRST CPU_TMS CPU_TDO CPU_TDI __3.3V __3.3V CPU_TCK CPU_FT_TDI CPU_FT_TDO CPU_FT_TMS CPU_FT_TRST CPU_FT_RST unnamed unnamed TXB0108
  XR110 GND unnamed R
  XR109 GND unnamed R
  XU6 GND GND GND _CPU_USB_JTAG_1.8V GND unnamed GND CPU_FT_TCK CPU_FT_TDI CPU_FT_TDO CPU_FT_TMS CPU_FT_XTIN __3.3V unnamed unnamed unnamed unnamed GND CPU_FT_TRST CPU_FT_RST CPU_FT_OE unnamed CPU_FT_XTOUT unnamed __3.3V unnamed unnamed unnamed GND unnamed _CPU_USB_JTAG_1.8V CPU_U2_RXD CPU_U2_TXD unnamed unnamed unnamed __3.3V unnamed unnamed unnamed unnamed GND unnamed _CPU_USB_JTAG_1.8V GND __3.3V GND unnamed unnamed unnamed unnamed __3.3V unnamed unnamed unnamed unnamed unnamed CPU_EEDATA CPU_EECLK CPU_EECS _CPU_USB_JTAG_1.8V CPU_USB_JTAG_DM CPU_USB_JTAG_DP unnamed FT2232H
  XC35 _CPU_USB_JTAG_1.8V GND C
  XFB7 unnamed __3.3V FILTER
  XC36 unnamed GND C
  XC38 unnamed GND C
  XC41 _CPU_USB_JTAG_1.8V GND C
  XC42 _CPU_USB_JTAG_1.8V GND C
  XC43 _CPU_USB_JTAG_1.8V GND C
  XC44 __3.3V GND C
  XC45 __3.3V GND C
  XC46 __3.3V GND C
  XC47 __3.3V GND C
  XR103 GND unnamed R
  XR104 __3.3V unnamed R
  XFB8 unnamed __3.3V FILTER
  XBT1 unnamed GND BATTERY
  XJP5 GND unnamed JUMPER
  XFB6 unnamed CPU_USB_DEBUG_VBUS FILTER
  XTR2 unnamed CPU_USB_JTAG_DP CPU_USB_JTAG_DM unnamed TRASF_UNIP
  XFB5 CPU_CHJ3 GND FILTER
  XC39 unnamed GND CAPAPOL
  XC37 unnamed GND CAPAPOL
  XJ3 unnamed unnamed unnamed GND GND CPU_CHJ3 CPU_CHJ3 CPU_CHJ3 CPU_CHJ3 CONN_9
  XR11 CPU_nTRST CPU_TRST R
  XR15 CPU_RESET CPU_RST R
  XFB9 GND unnamed FILTER
  XU8 CPU_CHJ3 CPU_USB_JTAG_DP CPU_USB_JTAG_DM unnamed PRTR5V0U2X
  XX1 CPU_RTCX2 unnamed unnamed CPU_RTCX1 CRYSTAL_4PIN_MINI_GND
  XFB10 unnamed __3.3VADC FILTER
  XD11 unnamed CPU_RESET DIODE
  XX2 CPU_XTAL1 GND CPU_XTAL2 GND SMD_SEALING_GLASS_CRYSTAL
  XX3 CPU_FT_XTOUT GND CPU_FT_XTIN GND SMD_SEALING_GLASS_CRYSTAL
  XC51 unnamed GND C
  XSW1 unnamed unnamed GND GND SW_PUSH
  XR58 CPU_PULS_0 unnamed R
  XR62 __3.3V unnamed R
  XC7 unnamed GND C
  XSW2 unnamed unnamed GND GND SW_PUSH
  XR59 CPU_PULS_1 unnamed R
  XR63 __3.3V unnamed R
  XC8 unnamed GND C
  XSW3 unnamed unnamed GND GND SW_PUSH
  XR60 CPU_PULS_2 unnamed R
  XR64 __3.3V unnamed R
  XC9 unnamed GND C
  XSW4 unnamed unnamed GND GND SW_PUSH
  XR61 CPU_PULS_3 unnamed R
  XR65 __3.3V unnamed R
  XC10 unnamed GND C
  XQ9 unnamed unnamed GND MOSFET_N
  XR82 CPU_LED1 unnamed R
  XR84 unnamed unnamed R
  XQ1 unnamed unnamed GND MOSFET_N
  XR66 CPU_LED0_B unnamed R
  XR68 unnamed unnamed R
  XQ3 unnamed unnamed GND MOSFET_N
  XR70 CPU_LED0_G unnamed R
  XR72 unnamed unnamed R
  XQ5 unnamed unnamed GND MOSFET_N
  XR74 CPU_LED0_R unnamed R
  XR76 unnamed unnamed R
  XQ4 unnamed unnamed GND MOSFET_N
  XR71 CPU_LED2 unnamed R
  XR73 unnamed unnamed R
  XLED1 unnamed unnamed unnamed _5V LED_ARBG
  XR12 CPU_LED0_G GND R
  XR14 CPU_LED0_R GND R
  XR10 CPU_LED0_B GND R
  XR18 CPU_LED1 GND R
  XR13 CPU_LED2 GND R
  XR19 CPU_LED3 GND R
  XR85 unnamed unnamed R
  XR83 CPU_LED3 unnamed R
  XQ10 unnamed unnamed GND MOSFET_N
  XD7 _5V unnamed LED
  XD9 _5V unnamed LED
  XD8 _5V unnamed LED
.ends \edu-ciaa-nxp

*--- Subcircuit Definitions ---
.subckt CONN_1 \1
* Stub for CONN_1
.ends

.subckt MAX3072 \1 \2 \3 \4 \5 \6 \7 \8
* Stub for MAX3072
.ends

.subckt C_MINI \1 \2
* Stub for C_MINI
.ends

.subckt R_MINI \1 \2
* Stub for R_MINI
.ends

.subckt ESD \1 \2
* Stub for ESD
.ends

.subckt \JUMPER-2 \1 \2
* Stub for \JUMPER-2
.ends

.subckt TB_1X3 \1 \2 \3
* Stub for TB_1X3
.ends

.subckt CP_MINI \1 \2
* Stub for CP_MINI
.ends

.subckt R \1 \2
* Stub for R
.ends

.subckt PRTR5V0U2X \1 \2 \3 \4
* Stub for PRTR5V0U2X
.ends

.subckt CAPAPOL \1 \2
* Stub for CAPAPOL
.ends

.subckt C \1 \2
* Stub for C
.ends

.subckt CONN_9 \1 \2 \3 \4 \5 \6 \7 \8 \9
* Stub for CONN_9
.ends

.subckt FILTER \1 \2
* Stub for FILTER
.ends

.subckt TRASF_UNIP \1 \2 \3 \4
* Stub for TRASF_UNIP
.ends

.subckt MIC2025 \1 \2 \3 \4 \5 \6 \7 \8
* Stub for MIC2025
.ends

.subckt THERMISTOR \1 \2
* Stub for THERMISTOR
.ends

.subckt CONN_20X2 \1 \10 \11 \12 \13 \14 \15 \16 \17 \18 \19 \2 \20 \21 \22 \23 \24 \25 \26 \27 \28 \29 \3 \30 \31 \32 \33 \34 \35 \36 \37 \38 \39 \4 \40 \5 \6 \7 \8 \9
* Stub for CONN_20X2
.ends

.subckt LED \1 \2
* Stub for LED
.ends

.subckt DIODESCH \1 \2
* Stub for DIODESCH
.ends

.subckt NCP1117ST15T3G \1 \2 \3 \4
* Stub for NCP1117ST15T3G
.ends

.subckt ZENER \1 \2
* Stub for ZENER
.ends

.subckt CONN_2 \1 \2
* Stub for CONN_2
.ends

.subckt SW_PUSH \1 \2 \3 \4
* Stub for SW_PUSH
.ends

.subckt LPC4337JBD144 \1 \10 \100 \101 \102 \103 \104 \105 \106 \107 \108 \109 \11 \110 \111 \112 \113 \114 \115 \116 \117 \118 \119 \12 \120 \121 \122 \123 \124 \125 \126 \127 \128 \129 \13 \130 \131 \132 \133 \134 \135 \136 \137 \138 \139 \14 \140 \141 \142 \143 \144 \15 \16 \17 \18 \19 \2 \20 \21 \22 \23 \24 \25 \26 \27 \28 \29 \3 \30 \31 \32 \33 \34 \35 \36 \37 \38 \39 \4 \40 \41 \42 \43 \44 \45 \46 \47 \48 \49 \5 \50 \51 \52 \53 \54 \55 \56 \57 \58 \59 \6 \60 \61 \62 \63 \64 \65 \66 \67 \68 \69 \7 \70 \71 \72 \73 \74 \75 \76 \77 \78 \79 \8 \80 \81 \82 \83 \84 \85 \86 \87 \88 \89 \9 \90 \91 \92 \93 \94 \95 \96 \97 \98 \99
* Stub for LPC4337JBD144
.ends

.subckt CONN_5X2 \1 \10 \2 \3 \4 \5 \6 \7 \8 \9
* Stub for CONN_5X2
.ends

.subckt \93C56 \1 \2 \3 \4 \5 \6 \7 \8
* Stub for \93C56
.ends

.subckt TXB0108 \1 \10 \11 \12 \13 \14 \15 \16 \17 \18 \19 \2 \20 \3 \4 \5 \6 \7 \8 \9
* Stub for TXB0108
.ends

.subckt FT2232H \1 \10 \11 \12 \13 \14 \15 \16 \17 \18 \19 \2 \20 \21 \22 \23 \24 \25 \26 \27 \28 \29 \3 \30 \31 \32 \33 \34 \35 \36 \37 \38 \39 \4 \40 \41 \42 \43 \44 \45 \46 \47 \48 \49 \5 \50 \51 \52 \53 \54 \55 \56 \57 \58 \59 \6 \60 \61 \62 \63 \64 \7 \8 \9
* Stub for FT2232H
.ends

.subckt BATTERY \1 \2
* Stub for BATTERY
.ends

.subckt JUMPER \1 \2
* Stub for JUMPER
.ends

.subckt CRYSTAL_4PIN_MINI_GND \1 \2 \3 \4
* Stub for CRYSTAL_4PIN_MINI_GND
.ends

.subckt DIODE \1 \2
* Stub for DIODE
.ends

.subckt SMD_SEALING_GLASS_CRYSTAL \1 \2 \3 \4
* Stub for SMD_SEALING_GLASS_CRYSTAL
.ends

.subckt MOSFET_N D G S
* Stub for MOSFET_N
.ends

.subckt LED_ARBG \1 \2 \3 \4
* Stub for LED_ARBG
.ends

