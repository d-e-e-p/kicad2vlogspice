//--- Top Level ---
module instance_array();



endmodule

//--- Cell Definitions ---
