* Spice Netlist (renamed)

*--- Top Level ---
.subckt edu-ciaa-nxp 
.ends edu-ciaa-nxp

