//--- Top Level ---
module div();



endmodule

//--- Cell Definitions ---
