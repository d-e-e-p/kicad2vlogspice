//--- Top Level ---
module ATMEGA328_Motor_Board();



endmodule

//--- Cell Definitions ---
