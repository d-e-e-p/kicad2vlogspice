* Spice Netlist (renamed)

*--- Top Level ---
.subckt instance_array 
.ends instance_array

