//--- Top Level ---
module \edu-ciaa-nxp ();



endmodule

//--- Cell Definitions ---
