//--- Top Level ---
module \A64-OlinuXino_Rev_H ();



endmodule

//--- Cell Definitions ---
