//--- Top Level ---
module HDMI2USB();



endmodule

//--- Cell Definitions ---
