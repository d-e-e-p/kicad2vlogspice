* Spice Netlist (renamed)

*--- Top Level ---
.subckt A64-OlinuXino_Rev_H AP_CK32KO AP_NMI_ AP_RESET_ GND GNDA IPS KEYADC NAND_Flash___eMMC__T_Card_and_Audio_HPOUTFB NAND_Flash___eMMC__T_Card_and_Audio_HPOUTL NAND_Flash___eMMC__T_Card_and_Audio_HPOUTR NAND_Flash___eMMC__T_Card_and_Audio_HP_DET NAND_Flash___eMMC__T_Card_and_Audio_LINEINL NAND_Flash___eMMC__T_Card_and_Audio_LINEINR NAND_Flash___eMMC__T_Card_and_Audio_LINEOUTL NAND_Flash___eMMC__T_Card_and_Audio_LINEOUTR NAND_Flash___eMMC__T_Card_and_Audio_MBIAS NAND_Flash___eMMC__T_Card_and_Audio_MICIN1N NAND_Flash___eMMC__T_Card_and_Audio_MICIN1P NAND_Flash___eMMC__T_Card_and_Audio_MICIN2N NAND_Flash___eMMC__T_Card_and_Audio_MICIN2P NAND_Flash___eMMC__T_Card_and_Audio_NAND0_ALE__SDC2_DS NAND_Flash___eMMC__T_Card_and_Audio_NAND0_DQ0__SDC2_D0 NAND_Flash___eMMC__T_Card_and_Audio_NAND0_DQ1__SDC2_D1 NAND_Flash___eMMC__T_Card_and_Audio_NAND0_DQ2__SDC2_D2 NAND_Flash___eMMC__T_Card_and_Audio_NAND0_DQ3__SDC2_D3 NAND_Flash___eMMC__T_Card_and_Audio_NAND0_DQ4__SDC2_D4 NAND_Flash___eMMC__T_Card_and_Audio_NAND0_DQ5__SDC2_D5 NAND_Flash___eMMC__T_Card_and_Audio_NAND0_DQ6__SDC2_D6 NAND_Flash___eMMC__T_Card_and_Audio_NAND0_DQ7__SDC2_D7 NAND_Flash___eMMC__T_Card_and_Audio_NAND0_DQS__SDC2_RST NAND_Flash___eMMC__T_Card_and_Audio_NAND0_RB0__SDC2_CMD NAND_Flash___eMMC__T_Card_and_Audio_NAND0_RE__SDC2_CLK NAND_Flash___eMMC__T_Card_and_Audio_SDC0_CLK NAND_Flash___eMMC__T_Card_and_Audio_SDC0_CMD NAND_Flash___eMMC__T_Card_and_Audio_SDC0_D0 NAND_Flash___eMMC__T_Card_and_Audio_SDC0_D1 NAND_Flash___eMMC__T_Card_and_Audio_SDC0_D2 NAND_Flash___eMMC__T_Card_and_Audio_SDC0_D3 NAND_Flash___eMMC__T_Card_and_Audio_SDC0_DET_ NAND_Flash___eMMC__T_Card_and_Audio_eMMC_CLK Net__3.3V_VCC_PE_2.8V1_Pad2_ Net__ANT1_Pad1_ Net__ANT2_Pad1_ Net__C105_Pad1_ Net__C105_Pad2_ Net__C107_Pad2_ Net__C125_Pad2_ Net__C135_Pad1_ Net__C143_Pad2_ Net__C149_Pad1_ Net__C151_Pad1_ Net__C174_Pad2_ Net__C177_Pad2_ Net__C181_Pad2_ Net__C182_Pad2_ Net__C183_Pad1_ Net__C184_Pad1_ Net__C185_Pad1_ Net__C187_Pad1_ Net__C188_Pad2_ Net__C192_Pad2_ Net__C196_Pad2_ Net__C198_Pad2_ Net__C199_Pad2_ Net__C200_Pad2_ Net__C204_Pad2_ Net__C207_Pad2_ Net__C211_Pad2_ Net__C212_Pad2_ Net__C213_Pad2_ Net__C218_Pad1_ Net__C37_Pad2_ Net__C42_Pad1_ Net__C45_Pad1_ Net__C48_Pad2_ Net__C51_Pad1_ Net__C52_Pad1_ Net__C54_Pad2_ Net__C55_Pad1_ Net__C57_Pad2_ Net__C58_Pad1_ Net__C59_Pad1_ Net__C60_Pad1_ Net__C61_Pad1_ Net__C61_Pad2_ Net__C62_Pad1_ Net__C63_Pad1_ Net__C64_Pad1_ Net__C65_Pad2_ Net__C66_Pad2_ Net__C68_Pad2_ Net__C74_Pad1_ Net__C75_Pad2_ Net__C86_Pad2_ Net__C87_Pad2_ Net__C88_Pad2_ Net__CHGLED1_Pad1_ Net__D2_Pad2_ Net__D3_Pad1_ Net__D4_Pad1_ Net__D4_Pad2_ Net__DBG_UART1_Pad1_ Net__FET1_Pad3_ Net__FET2_Pad1_ Net__FET3_Pad1_ Net__GPIO_LED1_Pad2_ Net__HDMI1_Pad14_ Net__HDMI1_Pad19_ Net__HEADPHONES_LINEOUT1_Pad1_ Net__HEADPHONES_LINEOUT1_Pad2_ Net__HEADPHONES_LINEOUT1_Pad3_ Net__HEADPHONES_LINEOUT1_Pad4_ Net__HEADPHONES_LINEOUT1_Pad5_ Net__HPHONEOUTL_LINEOUTL1_Pad2_ Net__HPHONEOUTR_LINEOUTR1_Pad2_ Net__HSIC1_Pad1_ Net__HSIC1_Pad2_ Net__HSIC1_Pad3_ Net__L14_Pad1_ Net__L15_Pad1_ Net__L17_Pad1_ Net__L18_Pad2_ Net__L19_Pad1_ Net__L20_Pad1_ Net__LINEINL_MICIN2_Pad2_ Net__LINEINR_MICIN1_Pad2_ Net__MICRO_SD1_Pad5_ Net__MIC_LINEIN1_Pad4_ Net__MIC_LINEIN1_Pad5_ Net__MIPI_DSI1_Pad16_ Net__MIPI_DSI1_Pad17_ Net__MIPI_DSI1_Pad19_ Net__MIPI_DSI1_Pad20_ Net__PWRLED1_Pad2_ Net__PWRON1_Pad1_ Net__R105_Pad2_ Net__R107_Pad1_ Net__R109_Pad2_ Net__R10_Pad1_ Net__R111_Pad2_ Net__R113_Pad2_ Net__R115_Pad1_ Net__R119_Pad1_ Net__R13_Pad1_ Net__R14_Pad1_ Net__R15_Pad1_ Net__R19_Pad1_ Net__R3_Pad2_ Net__R41_Pad2_ Net__R49_Pad2_ Net__R4_Pad2_ Net__R54_Pad1_ Net__R55_Pad1_ Net__R57_Pad1_ Net__R60_Pad1_ Net__R72_Pad1_ Net__R7_Pad2_ Net__R80_Pad2_ Net__R82_Pad1_ Net__R83_Pad1_ Net__R86_Pad1_ Net__R87_Pad1_ Net__R89_Pad1_ Net__R94_Pad1_ Net__R96_Pad1_ Net__R97_Pad1_ Net__R98_Pad1_ Net__R9_Pad1_ Net__RM15_Pad1.1_ Net__RM15_Pad2.1_ Net__RM15_Pad3.1_ Net__RM15_Pad4.1_ Net__RM1_Pad1.2_ Net__RM1_Pad2.2_ Net__RM1_Pad3.2_ Net__RM1_Pad4.2_ Net__T1_Pad3_ Net__U11_Pad10_ Net__U11_Pad11_ Net__U11_Pad21_ Net__U11_Pad23_ Net__U11_Pad29_ Net__U11_Pad30_ Net__U11_Pad32_ Net__U11_Pad35_ Net__U11_Pad37_ Net__U11_Pad38_ Net__U11_Pad39_ Net__U11_Pad3_ Net__U11_Pad40_ Net__U11_Pad4_ Net__U11_Pad5_ Net__U11_Pad8_ Net__U13_Pad6_ Net__U14_Pad23_ Net__U14_Pad24_ Net__U15_Pad13_ Net__U15_Pad43_ Net__U15_Pad47_ Net__U1_PadA13_ Net__U1_PadB10_ Net__U1_PadB13_ Net__U1_PadC14_ Net__U1_PadD14_ Net__U1_PadE16_ Net__U1_PadF16_ PC4 PC7 PH10 PH11 PL10 PL11 PL12 PL7 PL8 PL9 PMU_SCK PMU_SDA Power_Supply__Extensions_and_MiPi_DSI_1.8V_DVDD_CSI Power_Supply__Extensions_and_MiPi_DSI_2.8V_AVDD_CSI Power_Supply__Extensions_and_MiPi_DSI_3.3V_MIPI Power_Supply__Extensions_and_MiPi_DSI_DC5SET Power_Supply__Extensions_and_MiPi_DSI_DSI_CKN Power_Supply__Extensions_and_MiPi_DSI_DSI_CKP Power_Supply__Extensions_and_MiPi_DSI_DSI_D0N Power_Supply__Extensions_and_MiPi_DSI_DSI_D0P Power_Supply__Extensions_and_MiPi_DSI_DSI_D1N Power_Supply__Extensions_and_MiPi_DSI_DSI_D1P Power_Supply__Extensions_and_MiPi_DSI_DSI_D2N Power_Supply__Extensions_and_MiPi_DSI_DSI_D2P Power_Supply__Extensions_and_MiPi_DSI_DSI_D3N Power_Supply__Extensions_and_MiPi_DSI_DSI_D3P Power_Supply__Extensions_and_MiPi_DSI_MIPI_DSI_BKL Power_Supply__Extensions_and_MiPi_DSI_MIPI_DSI_EN Power_Supply__Extensions_and_MiPi_DSI_MIPI_DSI_RST Power_Supply__Extensions_and_MiPi_DSI_PB0 Power_Supply__Extensions_and_MiPi_DSI_PB1 Power_Supply__Extensions_and_MiPi_DSI_PB2 Power_Supply__Extensions_and_MiPi_DSI_PB3 Power_Supply__Extensions_and_MiPi_DSI_PB4 Power_Supply__Extensions_and_MiPi_DSI_PE0 Power_Supply__Extensions_and_MiPi_DSI_PE1 Power_Supply__Extensions_and_MiPi_DSI_PE10 Power_Supply__Extensions_and_MiPi_DSI_PE11 Power_Supply__Extensions_and_MiPi_DSI_PE12 Power_Supply__Extensions_and_MiPi_DSI_PE13 Power_Supply__Extensions_and_MiPi_DSI_PE14 Power_Supply__Extensions_and_MiPi_DSI_PE15 Power_Supply__Extensions_and_MiPi_DSI_PE16 Power_Supply__Extensions_and_MiPi_DSI_PE16__POWERON Power_Supply__Extensions_and_MiPi_DSI_PE17__GPIO_LED Power_Supply__Extensions_and_MiPi_DSI_PE2 Power_Supply__Extensions_and_MiPi_DSI_PE3 Power_Supply__Extensions_and_MiPi_DSI_PE4 Power_Supply__Extensions_and_MiPi_DSI_PE5 Power_Supply__Extensions_and_MiPi_DSI_PE6 Power_Supply__Extensions_and_MiPi_DSI_PE7 Power_Supply__Extensions_and_MiPi_DSI_PE8 Power_Supply__Extensions_and_MiPi_DSI_PE9 Power_Supply__Extensions_and_MiPi_DSI_UEXT_CLK Power_Supply__Extensions_and_MiPi_DSI_UEXT_CS Power_Supply__Extensions_and_MiPi_DSI_UEXT_MISO Power_Supply__Extensions_and_MiPi_DSI_UEXT_MOSI S0SA0 S0SA1 S0SA10 S0SA11 S0SA12 S0SA13 S0SA14 S0SA15 S0SA2 S0SA3 S0SA4 S0SA5 S0SA6 S0SA7 S0SA8 S0SA9 S0SBA0 S0SBA1 S0SBA2 S0SCAS S0SCKE0 S0SCKE1 S0SCK_N S0SCK_P S0SCS0 S0SCS1 S0SDQ0 S0SDQ1 S0SDQ10 S0SDQ11 S0SDQ12 S0SDQ13 S0SDQ14 S0SDQ15 S0SDQ16 S0SDQ17 S0SDQ18 S0SDQ19 S0SDQ2 S0SDQ20 S0SDQ21 S0SDQ22 S0SDQ23 S0SDQ24 S0SDQ25 S0SDQ26 S0SDQ27 S0SDQ28 S0SDQ29 S0SDQ3 S0SDQ30 S0SDQ31 S0SDQ4 S0SDQ5 S0SDQ6 S0SDQ7 S0SDQ8 S0SDQ9 S0SDQM0 S0SDQM1 S0SDQM2 S0SDQM3 S0SDQS0_N S0SDQS0_P S0SDQS1_N S0SDQS1_P S0SDQS2_N S0SDQS2_P S0SDQS3_N S0SDQS3_P S0SODT0 S0SODT1 S0SRAS S0SRST S0SVREF S0SWE SPI0_CLK SPI0_CS SPI0_MISO SPI0_MOSI TWI0_SCK TWI0_SDA TWI1_SCK TWI1_SDA UART3_RX UART3_TX UBOOT USB0_DRV USB0_D_N USB0_D_P USB1_DRV USB_HDMI_WiFi_BT_Ethernet_LCD_1.25_EXT USB_HDMI_WiFi_BT_Ethernet_LCD_AP_WAKE_BT USB_HDMI_WiFi_BT_Ethernet_LCD_BT_PCM_CLK USB_HDMI_WiFi_BT_Ethernet_LCD_BT_PCM_DIN USB_HDMI_WiFi_BT_Ethernet_LCD_BT_PCM_DOUT USB_HDMI_WiFi_BT_Ethernet_LCD_BT_PCM_SYNC USB_HDMI_WiFi_BT_Ethernet_LCD_BT_RST_N USB_HDMI_WiFi_BT_Ethernet_LCD_BT_UART_CTS USB_HDMI_WiFi_BT_Ethernet_LCD_BT_UART_RX USB_HDMI_WiFi_BT_Ethernet_LCD_BT_UART_TX USB_HDMI_WiFi_BT_Ethernet_LCD_BT_WAKE_AP USB_HDMI_WiFi_BT_Ethernet_LCD_EPHY_RST_ USB_HDMI_WiFi_BT_Ethernet_LCD_GCLKIN_LCD_VSYNC USB_HDMI_WiFi_BT_Ethernet_LCD_GMDC_LCD_PWM USB_HDMI_WiFi_BT_Ethernet_LCD_GMDIO_LCD_PWR USB_HDMI_WiFi_BT_Ethernet_LCD_GRXCK_LCD_D18 USB_HDMI_WiFi_BT_Ethernet_LCD_GRXCTL_LCD_D19 USB_HDMI_WiFi_BT_Ethernet_LCD_GRXD0_LCD_D15 USB_HDMI_WiFi_BT_Ethernet_LCD_GRXD1_LCD_D14 USB_HDMI_WiFi_BT_Ethernet_LCD_GRXD2_LCD_D13 USB_HDMI_WiFi_BT_Ethernet_LCD_GRXD3_LCD_D12 USB_HDMI_WiFi_BT_Ethernet_LCD_GTXCK_LCD_DE USB_HDMI_WiFi_BT_Ethernet_LCD_GTXCTL_LCD_HSYNC USB_HDMI_WiFi_BT_Ethernet_LCD_GTXD0_LCD_CLK USB_HDMI_WiFi_BT_Ethernet_LCD_GTXD1_LCD_D23 USB_HDMI_WiFi_BT_Ethernet_LCD_GTXD2_LCD_D22 USB_HDMI_WiFi_BT_Ethernet_LCD_GTXD3_LCD_D21 USB_HDMI_WiFi_BT_Ethernet_LCD_HCEC USB_HDMI_WiFi_BT_Ethernet_LCD_HHPD USB_HDMI_WiFi_BT_Ethernet_LCD_HSCL USB_HDMI_WiFi_BT_Ethernet_LCD_HSDA USB_HDMI_WiFi_BT_Ethernet_LCD_HTX0N USB_HDMI_WiFi_BT_Ethernet_LCD_HTX0P USB_HDMI_WiFi_BT_Ethernet_LCD_HTX1N USB_HDMI_WiFi_BT_Ethernet_LCD_HTX1P USB_HDMI_WiFi_BT_Ethernet_LCD_HTX2N USB_HDMI_WiFi_BT_Ethernet_LCD_HTX2P USB_HDMI_WiFi_BT_Ethernet_LCD_HTXCN USB_HDMI_WiFi_BT_Ethernet_LCD_HTXCP USB_HDMI_WiFi_BT_Ethernet_LCD_LCD_D10 USB_HDMI_WiFi_BT_Ethernet_LCD_LCD_D11 USB_HDMI_WiFi_BT_Ethernet_LCD_LCD_D2 USB_HDMI_WiFi_BT_Ethernet_LCD_LCD_D20 USB_HDMI_WiFi_BT_Ethernet_LCD_LCD_D3 USB_HDMI_WiFi_BT_Ethernet_LCD_LCD_D4 USB_HDMI_WiFi_BT_Ethernet_LCD_LCD_D5 USB_HDMI_WiFi_BT_Ethernet_LCD_LCD_D6 USB_HDMI_WiFi_BT_Ethernet_LCD_LCD_D7 USB_HDMI_WiFi_BT_Ethernet_LCD_MDI_0__ USB_HDMI_WiFi_BT_Ethernet_LCD_MDI_0___0 USB_HDMI_WiFi_BT_Ethernet_LCD_MDI_1__ USB_HDMI_WiFi_BT_Ethernet_LCD_MDI_1___0 USB_HDMI_WiFi_BT_Ethernet_LCD_MDI_2__ USB_HDMI_WiFi_BT_Ethernet_LCD_MDI_2___0 USB_HDMI_WiFi_BT_Ethernet_LCD_MDI_3__ USB_HDMI_WiFi_BT_Ethernet_LCD_MDI_3___0 USB_HDMI_WiFi_BT_Ethernet_LCD_PH7_CTP_INT USB_HDMI_WiFi_BT_Ethernet_LCD_PH8_CTP_RST USB_HDMI_WiFi_BT_Ethernet_LCD_PHYAD0 USB_HDMI_WiFi_BT_Ethernet_LCD_PHYAD1 USB_HDMI_WiFi_BT_Ethernet_LCD_USB0_ID USB_HDMI_WiFi_BT_Ethernet_LCD_USB0_VBUSDET USB_HDMI_WiFi_BT_Ethernet_LCD_USB1_DM USB_HDMI_WiFi_BT_Ethernet_LCD_USB1_DP USB_HDMI_WiFi_BT_Ethernet_LCD_VDD33 USB_HDMI_WiFi_BT_Ethernet_LCD_WL_PMU_EN USB_HDMI_WiFi_BT_Ethernet_LCD_WL_SDIO_CLK USB_HDMI_WiFi_BT_Ethernet_LCD_WL_SDIO_CMD USB_HDMI_WiFi_BT_Ethernet_LCD_WL_SDIO_D0 USB_HDMI_WiFi_BT_Ethernet_LCD_WL_SDIO_D1 USB_HDMI_WiFi_BT_Ethernet_LCD_WL_SDIO_D2 USB_HDMI_WiFi_BT_Ethernet_LCD_WL_SDIO_D3 USB_HDMI_WiFi_BT_Ethernet_LCD_WL_WAKE_AP VBAT VCC_PC VCC_PE VCC_PL VDDFB_CPUX VREF0_DDR3 _1.1V_CPUS _1.1V_CPUX _1.1V_SYS _1.2V_HSIC _1.5V _1.8V _3.0VA _3.0V_RTC _3.3V _3.3VD _3.3VWiFiIO _5V _5V_EXT _5V_USBOTG
  XC31 _1.5V GND C
  XC28 _1.5V GND C
  XC27 _1.5V GND C
  XC26 _1.5V GND C
  XC30 _1.5V GND C
  XC29 _1.5V GND C
  XR7 GND Net__R7_Pad2_ R
  XC22 GND S0SVREF C
  XR3 S0SCK_P Net__R3_Pad2_ R
  XR4 S0SCK_N Net__R4_Pad2_ R
  XR9 Net__R9_Pad1_ GND R
  XR13 Net__R13_Pad1_ GND R
  XR8 GND VREF0_DDR3 R
  XR5 VREF0_DDR3 _1.5V R
  XC11 _1.5V VREF0_DDR3 C
  XC23 VREF0_DDR3 GND C
  XC24 VREF0_DDR3 GND C
  XC12 _1.5V GND C
  XC13 _1.5V GND C
  XC14 _1.5V GND C
  XC15 _1.5V GND C
  XC16 _1.5V GND C
  XC1 _1.5V GND C
  XC2 _1.5V GND C
  XC3 _1.5V GND C
  XC4 _1.5V GND C
  XC5 _1.5V GND C
  XR12 GND S0SVREF R
  XR11 S0SVREF _1.5V R
  XC32 S0SVREF _1.5V C
  XC33 GND S0SVREF C
  XR10 Net__R10_Pad1_ GND R
  XR14 Net__R14_Pad1_ GND R
  XC25 VREF0_DDR3 GND C
  XC17 _1.5V GND C
  XC18 _1.5V GND C
  XC19 _1.5V GND C
  XC20 _1.5V GND C
  XC21 _1.5V GND C
  XC6 _1.5V GND C
  XC7 _1.5V GND C
  XC8 _1.5V GND C
  XC9 _1.5V GND C
  XC10 _1.5V GND C
  XR2 S0SCK_N S0SCK_P R
  XR1 S0SRST _1.5V R
  XR6 VREF0_DDR3 S0SVREF R
  XU2 _1.5V S0SDQ15 S0SDQ12 S0SDQ8 _1.5V GND GND _1.5V GND S0SDQS1_N S0SDQ10 GND _1.5V S0SDQ13 S0SDQ14 S0SDQS1_P S0SDQ9 _1.5V GND _1.5V S0SDQM1 S0SDQ11 GND _1.5V GND GND S0SDQ4 S0SDQM0 GND _1.5V _1.5V S0SDQ2 S0SDQS0_P S0SDQ0 S0SDQ7 GND GND S0SDQ1 S0SDQS0_N _1.5V GND GND VREF0_DDR3 _1.5V S0SDQ5 S0SDQ3 S0SDQ6 _1.5V S0SODT1 GND S0SRAS S0SCK_P GND S0SCKE1 S0SODT0 _1.5V S0SCAS S0SCK_N _1.5V S0SCKE0 S0SCS1 S0SCS0 S0SWE S0SA10 Net__R9_Pad1_ Net__R13_Pad1_ GND S0SBA0 S0SBA2 S0SA15 VREF0_DDR3 GND _1.5V S0SA3 S0SA0 S0SA12 S0SBA1 _1.5V GND S0SA5 S0SA2 S0SA1 S0SA4 GND _1.5V S0SA7 S0SA9 S0SA11 S0SA6 _1.5V GND S0SRST S0SA13 S0SA14 S0SA8 GND H5TQ2G63BFR_MEM4G16D3EABG-125--H5TC8G63AMR-PBA_K4B8G1646Q-MYK0(FBGA-96_512MX16_DDR3-1600_11-11-11)
  XU3 _1.5V S0SDQ30 S0SDQ28 S0SDQ24 _1.5V GND GND _1.5V GND S0SDQS3_N S0SDQ27 GND _1.5V S0SDQ31 S0SDQ29 S0SDQS3_P S0SDQ25 _1.5V GND _1.5V S0SDQM3 S0SDQ26 GND _1.5V GND GND S0SDQ22 S0SDQM2 GND _1.5V _1.5V S0SDQ21 S0SDQS2_P S0SDQ16 S0SDQ19 GND GND S0SDQ23 S0SDQS2_N _1.5V GND GND VREF0_DDR3 _1.5V S0SDQ20 S0SDQ18 S0SDQ17 _1.5V S0SODT1 GND S0SRAS S0SCK_P GND S0SCKE1 S0SODT0 _1.5V S0SCAS S0SCK_N _1.5V S0SCKE0 S0SCS1 S0SCS0 S0SWE S0SA10 Net__R10_Pad1_ Net__R14_Pad1_ GND S0SBA0 S0SBA2 S0SA15 VREF0_DDR3 GND _1.5V S0SA3 S0SA0 S0SA12 S0SBA1 _1.5V GND S0SA5 S0SA2 S0SA1 S0SA4 GND _1.5V S0SA7 S0SA9 S0SA11 S0SA6 _1.5V GND S0SRST S0SA13 S0SA14 S0SA8 GND H5TQ2G63BFR_MEM4G16D3EABG-125--H5TC8G63AMR-PBA_K4B8G1646Q-MYK0(FBGA-96_512MX16_DDR3-1600_11-11-11)
  XU1 GND GNDA Net__U1_PadA13_ NAND_Flash___eMMC__T_Card_and_Audio_LINEINR KEYADC NAND_Flash___eMMC__T_Card_and_Audio_MICIN2N USB_HDMI_WiFi_BT_Ethernet_LCD_WL_PMU_EN S0SDQ22 USB_HDMI_WiFi_BT_Ethernet_LCD_BT_RST_N USB0_D_P GND S0SDQ26 S0SDQ27 S0SDQ28 S0SDQ29 _1.1V_CPUX TWI0_SDA Net__R97_Pad1_ Net__R98_Pad1_ USB_HDMI_WiFi_BT_Ethernet_LCD_GRXD2_LCD_D13 USB_HDMI_WiFi_BT_Ethernet_LCD_LCD_D5 USB_HDMI_WiFi_BT_Ethernet_LCD_LCD_D7 USB_HDMI_WiFi_BT_Ethernet_LCD_LCD_D11 USB_HDMI_WiFi_BT_Ethernet_LCD_LCD_D3 Power_Supply__Extensions_and_MiPi_DSI_PE0 Power_Supply__Extensions_and_MiPi_DSI_PE4 USB_HDMI_WiFi_BT_Ethernet_LCD_LCD_D2 Power_Supply__Extensions_and_MiPi_DSI_PE3 Power_Supply__Extensions_and_MiPi_DSI_PE2 _1.1V_CPUX PH11 Power_Supply__Extensions_and_MiPi_DSI_MIPI_DSI_RST Power_Supply__Extensions_and_MiPi_DSI_PB3 USB_HDMI_WiFi_BT_Ethernet_LCD_USB0_ID TWI1_SDA NAND_Flash___eMMC__T_Card_and_Audio_SDC0_D1 Net__R72_Pad1_ Net__R19_Pad1_ Net__RM1_Pad2.2_ Net__RM1_Pad4.2_ USB_HDMI_WiFi_BT_Ethernet_LCD_LCD_D20 USB_HDMI_WiFi_BT_Ethernet_LCD_GRXCTL_LCD_D19 USB_HDMI_WiFi_BT_Ethernet_LCD_BT_UART_RX USB_HDMI_WiFi_BT_Ethernet_LCD_BT_PCM_CLK USB_HDMI_WiFi_BT_Ethernet_LCD_BT_PCM_SYNC _1.1V_CPUX Power_Supply__Extensions_and_MiPi_DSI_PE12 Power_Supply__Extensions_and_MiPi_DSI_PE16 Power_Supply__Extensions_and_MiPi_DSI_PE10 Power_Supply__Extensions_and_MiPi_DSI_PE1 USB_HDMI_WiFi_BT_Ethernet_LCD_USB0_VBUSDET UART3_TX NAND_Flash___eMMC__T_Card_and_Audio_SDC0_D3 Power_Supply__Extensions_and_MiPi_DSI_PB1 NAND_Flash___eMMC__T_Card_and_Audio_SDC0_DET_ NAND_Flash___eMMC__T_Card_and_Audio_SDC0_D2 _1.1V_CPUX USB_HDMI_WiFi_BT_Ethernet_LCD_GMDIO_LCD_PWR USB_HDMI_WiFi_BT_Ethernet_LCD_GCLKIN_LCD_VSYNC Net__RM1_Pad1.2_ Net__RM1_Pad3.2_ USB_HDMI_WiFi_BT_Ethernet_LCD_GRXCK_LCD_D18 USB_HDMI_WiFi_BT_Ethernet_LCD_BT_UART_CTS USB_HDMI_WiFi_BT_Ethernet_LCD_BT_PCM_DIN _1.1V_CPUX Power_Supply__Extensions_and_MiPi_DSI_PE14 Power_Supply__Extensions_and_MiPi_DSI_PE8 GND TWI1_SCK USB_HDMI_WiFi_BT_Ethernet_LCD_PH7_CTP_INT UART3_RX NAND_Flash___eMMC__T_Card_and_Audio_SDC0_CLK S0SDQ20 Net__U1_PadB10_ Net__C59_Pad1_ Net__C55_Pad1_ Net__U1_PadB13_ NAND_Flash___eMMC__T_Card_and_Audio_LINEINL NAND_Flash___eMMC__T_Card_and_Audio_MICIN1P NAND_Flash___eMMC__T_Card_and_Audio_MICIN1N NAND_Flash___eMMC__T_Card_and_Audio_MICIN2P AP_CK32KO Net__C183_Pad1_ S0SDQ21 USB_HDMI_WiFi_BT_Ethernet_LCD_AP_WAKE_BT PL8 USB0_D_N USB_HDMI_WiFi_BT_Ethernet_LCD_USB1_DP S0SDQ23 S0SDQ25 S0SDQS3_N S0SDQS3_P S0SDQM3 S0SDQ30 S0SDQ31 NAND_Flash___eMMC__T_Card_and_Audio_HPOUTFB Net__C51_Pad1_ NAND_Flash___eMMC__T_Card_and_Audio_HPOUTR NAND_Flash___eMMC__T_Card_and_Audio_HPOUTL Net__U1_PadC14_ NAND_Flash___eMMC__T_Card_and_Audio_LINEOUTR PMU_SDA Net__C184_Pad1_ PL7 S0SDQM2 PL11 USB_HDMI_WiFi_BT_Ethernet_LCD_USB1_DM GND S0SA9 S0SDQ24 S0SBA2 GND S0SWE S0SCAS S0SDQS2_N S0SRST NAND_Flash___eMMC__T_Card_and_Audio_HP_DET Net__C63_Pad1_ Net__U1_PadD14_ NAND_Flash___eMMC__T_Card_and_Audio_LINEOUTL PMU_SCK USB_HDMI_WiFi_BT_Ethernet_LCD_BT_WAKE_AP S0SDQS2_P PL9 PL10 PL12 USB_HDMI_WiFi_BT_Ethernet_LCD_HTX2P S0SA8 S0SODT0 GND S0SBA0 S0SDQ19 Net__C61_Pad2_ Net__C61_Pad1_ _1.8V NAND_Flash___eMMC__T_Card_and_Audio_MBIAS Net__U1_PadE16_ AP_RESET_ USB_HDMI_WiFi_BT_Ethernet_LCD_WL_WAKE_AP S0SDQ18 USB_HDMI_WiFi_BT_Ethernet_LCD_HSDA USB_HDMI_WiFi_BT_Ethernet_LCD_HHPD USB_HDMI_WiFi_BT_Ethernet_LCD_HTX2N USB_HDMI_WiFi_BT_Ethernet_LCD_HTX1P S0SDQ16 S0SA7 S0SCS0 S0SODT1 S0SA13 Net__C54_Pad2_ Net__U1_PadF16_ UBOOT S0SDQ17 USB_HDMI_WiFi_BT_Ethernet_LCD_HCEC USB_HDMI_WiFi_BT_Ethernet_LCD_HTX1N S0SA6 S0SRAS S0SDQ1 GND Net__C54_Pad2_ _3.0VA Net__C192_Pad2_ AP_NMI_ Net__HSIC1_Pad3_ Net__R3_Pad2_ NAND_Flash___eMMC__T_Card_and_Audio_NAND0_RE__SDC2_CLK USB_HDMI_WiFi_BT_Ethernet_LCD_HSCL USB_HDMI_WiFi_BT_Ethernet_LCD_HTX0P USB_HDMI_WiFi_BT_Ethernet_LCD_HTX0N Net__R4_Pad2_ S0SA5 S0SVREF GND _1.5V _1.5V _1.5V S0SDQ5 GND Net__R96_Pad1_ _1.1V_CPUS _3.0V_RTC Net__HSIC1_Pad2_ S0SDQ4 NAND_Flash___eMMC__T_Card_and_Audio_NAND0_DQ3__SDC2_D3 USB_HDMI_WiFi_BT_Ethernet_LCD_HTXCP USB_HDMI_WiFi_BT_Ethernet_LCD_HTXCN S0SDQ2 GND S0SCS1 S0SCKE1 GND GND _1.1V_SYS _1.1V_SYS GND GND VCC_PL S0SDQM0 NAND_Flash___eMMC__T_Card_and_Audio_NAND0_DQ6__SDC2_D6 S0SCKE0 _1.5V GND S0SDQ3 GND GND GND GND _1.1V_SYS _1.2V_HSIC NAND_Flash___eMMC__T_Card_and_Audio_NAND0_ALE__SDC2_DS NAND_Flash___eMMC__T_Card_and_Audio_NAND0_RB0__SDC2_CMD S0SDQS0_N NAND_Flash___eMMC__T_Card_and_Audio_NAND0_DQ2__SDC2_D2 Net__C187_Pad1_ Net__R94_Pad1_ S0SDQS0_P S0SA14 S0SA12 _1.5V _1.5V GND GND S0SDQ6 GND GND GND _1.1V_SYS _1.1V_SYS GND _3.3V NAND_Flash___eMMC__T_Card_and_Audio_NAND0_DQ1__SDC2_D1 S0SDQ7 NAND_Flash___eMMC__T_Card_and_Audio_NAND0_DQ5__SDC2_D5 Power_Supply__Extensions_and_MiPi_DSI_DSI_D3N Power_Supply__Extensions_and_MiPi_DSI_DSI_D3P S0SDQ0 GND GND _1.5V _1.5V _1.5V GND GND GND GND _1.1V_SYS _1.1V_SYS GND _3.3VD S0SDQ15 NAND_Flash___eMMC__T_Card_and_Audio_NAND0_DQ0__SDC2_D0 Power_Supply__Extensions_and_MiPi_DSI_DSI_D2P GND S0SA10 GND GND S0SDQ14 GND GND GND GND _1.1V_SYS GND _3.0VA _3.3V _3.3V S0SDQ13 NAND_Flash___eMMC__T_Card_and_Audio_NAND0_DQS__SDC2_RST Power_Supply__Extensions_and_MiPi_DSI_DSI_D2N Power_Supply__Extensions_and_MiPi_DSI_DSI_CKP S0SDQ12 GND S0SA2 S0SA3 _1.5V _1.5V GND S0SDQS1_P GND GND GND GND _1.1V_SYS Net__C188_Pad2_ NAND_Flash___eMMC__T_Card_and_Audio_NAND0_DQ4__SDC2_D4 SPI0_CS S0SDQS1_N SPI0_CLK Power_Supply__Extensions_and_MiPi_DSI_DSI_D1P Power_Supply__Extensions_and_MiPi_DSI_DSI_CKN S0SDQM1 S0SA0 S0SA4 GND GND GND GND GND GND _1.1V_SYS _1.1V_SYS GND VCC_PC S0SDQ11 NAND_Flash___eMMC__T_Card_and_Audio_NAND0_DQ7__SDC2_D7 Power_Supply__Extensions_and_MiPi_DSI_DSI_D1N S0SBA1 S0SA1 GND GND GND GND GND S0SDQ10 GND GND GND GND _3.3V _1.1V_SYS _3.3VWiFiIO PC7 S0SDQ9 PC4 SPI0_MOSI Power_Supply__Extensions_and_MiPi_DSI_DSI_D0P Power_Supply__Extensions_and_MiPi_DSI_DSI_D0N S0SDQ8 S0SA15 VDDFB_CPUX GND GND Net__R7_Pad2_ GND GND _3.3V _3.3V Net__3.3V_VCC_PE_2.8V1_Pad2_ USB_HDMI_WiFi_BT_Ethernet_LCD_WL_SDIO_D0 GND USB_HDMI_WiFi_BT_Ethernet_LCD_WL_SDIO_CMD USB1_DRV USB_HDMI_WiFi_BT_Ethernet_LCD_BT_PCM_DOUT USB_HDMI_WiFi_BT_Ethernet_LCD_BT_UART_TX S0SA11 GND _1.1V_CPUX GND GND GND Net__DBG_UART1_Pad1_ GND USB_HDMI_WiFi_BT_Ethernet_LCD_GRXD3_LCD_D12 USB_HDMI_WiFi_BT_Ethernet_LCD_LCD_D6 _1.1V_CPUX USB_HDMI_WiFi_BT_Ethernet_LCD_WL_SDIO_CLK USB_HDMI_WiFi_BT_Ethernet_LCD_WL_SDIO_D1 _1.1V_CPUX _1.1V_CPUX _1.1V_CPUX _1.1V_CPUX GND Power_Supply__Extensions_and_MiPi_DSI_PB0 _1.1V_CPUX Power_Supply__Extensions_and_MiPi_DSI_PB2 TWI0_SCK NAND_Flash___eMMC__T_Card_and_Audio_SDC0_D0 USB_HDMI_WiFi_BT_Ethernet_LCD_GRXD1_LCD_D14 Power_Supply__Extensions_and_MiPi_DSI_PE5 USB_HDMI_WiFi_BT_Ethernet_LCD_LCD_D4 Power_Supply__Extensions_and_MiPi_DSI_PE6 Power_Supply__Extensions_and_MiPi_DSI_PE11 Power_Supply__Extensions_and_MiPi_DSI_PE17__GPIO_LED USB_HDMI_WiFi_BT_Ethernet_LCD_WL_SDIO_D3 _1.1V_CPUX _1.1V_CPUX _1.1V_CPUX Power_Supply__Extensions_and_MiPi_DSI_PB4 Power_Supply__Extensions_and_MiPi_DSI_MIPI_DSI_BKL NAND_Flash___eMMC__T_Card_and_Audio_SDC0_CMD USB_HDMI_WiFi_BT_Ethernet_LCD_PH8_CTP_RST USB_HDMI_WiFi_BT_Ethernet_LCD_LCD_D10 USB_HDMI_WiFi_BT_Ethernet_LCD_GMDC_LCD_PWM USB_HDMI_WiFi_BT_Ethernet_LCD_EPHY_RST_ USB_HDMI_WiFi_BT_Ethernet_LCD_GRXD0_LCD_D15 Power_Supply__Extensions_and_MiPi_DSI_PE9 Power_Supply__Extensions_and_MiPi_DSI_PE7 _1.1V_CPUX USB_HDMI_WiFi_BT_Ethernet_LCD_WL_SDIO_D2 Power_Supply__Extensions_and_MiPi_DSI_PE13 Power_Supply__Extensions_and_MiPi_DSI_PE15 _1.1V_CPUX _1.1V_CPUX Power_Supply__Extensions_and_MiPi_DSI_MIPI_DSI_EN Net__D4_Pad2_ PH10 AllWinner-A64(FBGA396)
  XC37 GND Net__C37_Pad2_ C
  XC38 GND Net__C37_Pad2_ C
  XC36 GND VCC_PC C
  XC35 GND VCC_PC C
  XC43 Net__C42_Pad1_ GND C
  XC44 Net__C42_Pad1_ GND C
  XL1 _3.3V Net__C42_Pad1_ L
  XC42 Net__C42_Pad1_ GND C
  XR21 NAND_Flash___eMMC__T_Card_and_Audio_NAND0_RB0__SDC2_CMD VCC_PC R
  XR23 NAND_Flash___eMMC__T_Card_and_Audio_NAND0_DQS__SDC2_RST VCC_PC R
  XC34 GND VCC_PC C
  XMICRO_SD1 NAND_Flash___eMMC__T_Card_and_Audio_SDC0_D2 GND GND GND GND NAND_Flash___eMMC__T_Card_and_Audio_SDC0_D3 NAND_Flash___eMMC__T_Card_and_Audio_SDC0_CMD Net__C64_Pad1_ Net__MICRO_SD1_Pad5_ GND NAND_Flash___eMMC__T_Card_and_Audio_SDC0_D0 NAND_Flash___eMMC__T_Card_and_Audio_SDC0_D1 NAND_Flash___eMMC__T_Card_and_Audio_SDC0_DET_ MICRO_SD(TFC-WPAPR-08)
  XR33 Net__MICRO_SD1_Pad5_ NAND_Flash___eMMC__T_Card_and_Audio_SDC0_CLK R
  XC64 Net__C64_Pad1_ GND C
  XL2 _3.3V Net__C64_Pad1_ L
  XRM7 _3.3V NAND_Flash___eMMC__T_Card_and_Audio_SDC0_D0 _3.3V NAND_Flash___eMMC__T_Card_and_Audio_SDC0_D1 _3.3V NAND_Flash___eMMC__T_Card_and_Audio_SDC0_DET_ _3.3V NAND_Flash___eMMC__T_Card_and_Audio_SDC0_D2 RA1206_(4x0603)_4B8_Smashed
  XR31 NAND_Flash___eMMC__T_Card_and_Audio_SDC0_CMD _3.3V R
  XR30 NAND_Flash___eMMC__T_Card_and_Audio_SDC0_D3 _3.3V R
  XC46 _3.0VA GNDA C
  XC49 _3.0VA GNDA C
  XC51 Net__C51_Pad1_ GNDA C
  XC53 Net__C51_Pad1_ GNDA C
  XC55 Net__C55_Pad1_ GNDA C
  XR27 Net__C59_Pad1_ GNDA R
  XC59 Net__C59_Pad1_ GNDA C
  XC63 Net__C63_Pad1_ GNDA C
  XMIC_LINEIN1 Net__LINEINL_MICIN2_Pad2_ GNDA Net__LINEINR_MICIN1_Pad2_ Net__MIC_LINEIN1_Pad4_ Net__MIC_LINEIN1_Pad5_ AUDIO_JACK(SCJ325P00XG0B02G)
  XC48 GNDA Net__C48_Pad2_ C
  XC62 Net__C62_Pad1_ GNDA C
  XC52 Net__C52_Pad1_ NAND_Flash___eMMC__T_Card_and_Audio_MICIN1P C
  XC60 Net__C60_Pad1_ NAND_Flash___eMMC__T_Card_and_Audio_MICIN2P C
  XR26 Net__C60_Pad1_ Net__C57_Pad2_ R
  XR25 Net__C57_Pad2_ NAND_Flash___eMMC__T_Card_and_Audio_MBIAS R
  XC57 GNDA Net__C57_Pad2_ C
  XR29 Net__C52_Pad1_ Net__C57_Pad2_ R
  XHEADPHONES_LINEOUT1 Net__HEADPHONES_LINEOUT1_Pad1_ Net__HEADPHONES_LINEOUT1_Pad2_ Net__HEADPHONES_LINEOUT1_Pad3_ Net__HEADPHONES_LINEOUT1_Pad4_ Net__HEADPHONES_LINEOUT1_Pad5_ AUDIO_JACK(SCJ325P00XG0B02G)
  XL3 Net__HPHONEOUTR_LINEOUTR1_Pad2_ Net__HEADPHONES_LINEOUT1_Pad3_ L
  XL4 NAND_Flash___eMMC__T_Card_and_Audio_HPOUTFB Net__HEADPHONES_LINEOUT1_Pad2_ L
  XL5 Net__HPHONEOUTL_LINEOUTL1_Pad2_ Net__HEADPHONES_LINEOUT1_Pad1_ L
  XC65 GNDA Net__C65_Pad2_ C
  XC66 GNDA Net__C66_Pad2_ C
  XR35 GNDA NAND_Flash___eMMC__T_Card_and_Audio_HPOUTR R
  XR32 Net__HEADPHONES_LINEOUT1_Pad4_ _3.0VA R
  XR34 GNDA NAND_Flash___eMMC__T_Card_and_Audio_HPOUTFB R
  XC61 Net__C61_Pad1_ Net__C61_Pad2_ C
  XC54 GNDA Net__C54_Pad2_ C
  XC56 GNDA Net__C54_Pad2_ C
  XC50 GNDA _1.8V C
  XC47 GNDA _1.8V C
  XR36 GND GNDA R
  XU12 SPI0_CS SPI0_MISO Net__R55_Pad1_ GND SPI0_MOSI SPI0_CLK Net__R57_Pad1_ _3.3V W25Q16BV
  XC81 GND _3.3V C
  XR57 Net__R57_Pad1_ _3.3V R
  XR56 Net__R55_Pad1_ _3.3V R
  XR55 Net__R55_Pad1_ GND R
  XR53 SPI0_CS _3.3V R
  XLINEINR_MICIN1 Net__C52_Pad1_ Net__LINEINR_MICIN1_Pad2_ Net__C45_Pad1_ SJ2W_Closed(1-2)
  XLINEINL_MICIN2 Net__C60_Pad1_ Net__LINEINL_MICIN2_Pad2_ Net__C58_Pad1_ SJ2W_Closed(1-2)
  XR59 Net__HEADPHONES_LINEOUT1_Pad4_ NAND_Flash___eMMC__T_Card_and_Audio_HP_DET R
  XR63 Net__C65_Pad2_ NAND_Flash___eMMC__T_Card_and_Audio_HPOUTL R
  XR64 Net__C66_Pad2_ NAND_Flash___eMMC__T_Card_and_Audio_HPOUTR R
  XHPHONEOUTR_LINEOUTR1 NAND_Flash___eMMC__T_Card_and_Audio_HPOUTR Net__HPHONEOUTR_LINEOUTR1_Pad2_ Net__C86_Pad2_ SJ2W_Closed(1-2)
  XHPHONEOUTL_LINEOUTL1 NAND_Flash___eMMC__T_Card_and_Audio_HPOUTL Net__HPHONEOUTL_LINEOUTL1_Pad2_ Net__C87_Pad2_ SJ2W_Closed(1-2)
  XC45 Net__C45_Pad1_ NAND_Flash___eMMC__T_Card_and_Audio_LINEINR C
  XC58 Net__C58_Pad1_ NAND_Flash___eMMC__T_Card_and_Audio_LINEINL C
  XC82 Net__C48_Pad2_ NAND_Flash___eMMC__T_Card_and_Audio_MICIN1N C
  XC83 Net__C62_Pad1_ NAND_Flash___eMMC__T_Card_and_Audio_MICIN2N C
  XC84 Net__C52_Pad1_ Net__C48_Pad2_ C
  XC85 Net__C60_Pad1_ Net__C62_Pad1_ C
  XC86 NAND_Flash___eMMC__T_Card_and_Audio_LINEOUTR Net__C86_Pad2_ C
  XC87 NAND_Flash___eMMC__T_Card_and_Audio_LINEOUTL Net__C87_Pad2_ C
  XGNDA1 GNDA TESTPAD
  XMounting_hole1 GND Mounting_hole
  XMounting_hole2 GND Mounting_hole
  XMounting_hole3 GND Mounting_hole
  XU5 NAND_Flash___eMMC__T_Card_and_Audio_NAND0_DQ0__SDC2_D0 NAND_Flash___eMMC__T_Card_and_Audio_NAND0_DQ1__SDC2_D1 NAND_Flash___eMMC__T_Card_and_Audio_NAND0_DQ2__SDC2_D2 GND NAND_Flash___eMMC__T_Card_and_Audio_NAND0_DQ3__SDC2_D3 NAND_Flash___eMMC__T_Card_and_Audio_NAND0_DQ4__SDC2_D4 NAND_Flash___eMMC__T_Card_and_Audio_NAND0_DQ5__SDC2_D5 NAND_Flash___eMMC__T_Card_and_Audio_NAND0_DQ6__SDC2_D6 NAND_Flash___eMMC__T_Card_and_Audio_NAND0_DQ7__SDC2_D7 Net__C37_Pad2_ GND VCC_PC Net__C42_Pad1_ GND Net__C42_Pad1_ GND GND Net__R15_Pad1_ Net__C42_Pad1_ GND NAND_Flash___eMMC__T_Card_and_Audio_NAND0_DQS__SDC2_RST GND Net__C42_Pad1_ VCC_PC NAND_Flash___eMMC__T_Card_and_Audio_NAND0_RB0__SDC2_CMD NAND_Flash___eMMC__T_Card_and_Audio_eMMC_CLK GND VCC_PC GND VCC_PC GND VCC_PC GND KLMAG2GEND-B031(FBGA153)
  XR67 NAND_Flash___eMMC__T_Card_and_Audio_NAND0_DQ0__SDC2_D0 VCC_PC R
  XWP_Enable1 GND Net__R55_Pad1_ SJ
  XR68 NAND_Flash___eMMC__T_Card_and_Audio_eMMC_CLK NAND_Flash___eMMC__T_Card_and_Audio_NAND0_RE__SDC2_CLK R
  XC94 NAND_Flash___eMMC__T_Card_and_Audio_eMMC_CLK GND C
  XR66 SPI0_MISO NAND_Flash___eMMC__T_Card_and_Audio_NAND0_ALE__SDC2_DS R
  XR62 NAND_Flash___eMMC__T_Card_and_Audio_NAND0_ALE__SDC2_DS GND R
  XR15 Net__R15_Pad1_ NAND_Flash___eMMC__T_Card_and_Audio_NAND0_ALE__SDC2_DS R
  XHDMI1 GND GND GND GND USB_HDMI_WiFi_BT_Ethernet_LCD_HTX2P USB_HDMI_WiFi_BT_Ethernet_LCD_HTXCP GND USB_HDMI_WiFi_BT_Ethernet_LCD_HTXCN Net__FET1_Pad3_ Net__HDMI1_Pad14_ USB_HDMI_WiFi_BT_Ethernet_LCD_HSCL USB_HDMI_WiFi_BT_Ethernet_LCD_HSDA GND Net__D3_Pad1_ Net__HDMI1_Pad19_ GND USB_HDMI_WiFi_BT_Ethernet_LCD_HTX2N USB_HDMI_WiFi_BT_Ethernet_LCD_HTX1P GND USB_HDMI_WiFi_BT_Ethernet_LCD_HTX1N USB_HDMI_WiFi_BT_Ethernet_LCD_HTX0P GND USB_HDMI_WiFi_BT_Ethernet_LCD_HTX0N HDMI-SWM-19
  XU7 USB_HDMI_WiFi_BT_Ethernet_LCD_HTX2P USB_HDMI_WiFi_BT_Ethernet_LCD_HTX2P USB_HDMI_WiFi_BT_Ethernet_LCD_HTX2N GND USB_HDMI_WiFi_BT_Ethernet_LCD_HTX1P USB_HDMI_WiFi_BT_Ethernet_LCD_HTX1N USB_HDMI_WiFi_BT_Ethernet_LCD_HTX1N USB_HDMI_WiFi_BT_Ethernet_LCD_HTX1P GND USB_HDMI_WiFi_BT_Ethernet_LCD_HTX2N RCLAMP0524P
  XU8 USB_HDMI_WiFi_BT_Ethernet_LCD_HTX0P USB_HDMI_WiFi_BT_Ethernet_LCD_HTX0P USB_HDMI_WiFi_BT_Ethernet_LCD_HTX0N GND USB_HDMI_WiFi_BT_Ethernet_LCD_HTXCP USB_HDMI_WiFi_BT_Ethernet_LCD_HTXCN USB_HDMI_WiFi_BT_Ethernet_LCD_HTXCN USB_HDMI_WiFi_BT_Ethernet_LCD_HTXCP GND USB_HDMI_WiFi_BT_Ethernet_LCD_HTX0N RCLAMP0524P
  XU10 USB_HDMI_WiFi_BT_Ethernet_LCD_HCEC USB_HDMI_WiFi_BT_Ethernet_LCD_HCEC USB_HDMI_WiFi_BT_Ethernet_LCD_HSCL GND USB_HDMI_WiFi_BT_Ethernet_LCD_HSDA USB_HDMI_WiFi_BT_Ethernet_LCD_HHPD USB_HDMI_WiFi_BT_Ethernet_LCD_HHPD USB_HDMI_WiFi_BT_Ethernet_LCD_HSDA GND USB_HDMI_WiFi_BT_Ethernet_LCD_HSCL RCLAMP0524P
  XR51 USB_HDMI_WiFi_BT_Ethernet_LCD_HHPD Net__HDMI1_Pad19_ R
  XR52 USB_HDMI_WiFi_BT_Ethernet_LCD_HHPD GND R
  XFET1 _3.3VD USB_HDMI_WiFi_BT_Ethernet_LCD_HCEC Net__FET1_Pad3_ N-MOS+DIOD_Small
  XR46 _3.3VD USB_HDMI_WiFi_BT_Ethernet_LCD_HCEC R
  XR50 _5V USB_HDMI_WiFi_BT_Ethernet_LCD_HSDA R
  XR47 _5V USB_HDMI_WiFi_BT_Ethernet_LCD_HSCL R
  XR39 USB_HDMI_WiFi_BT_Ethernet_LCD_HTX2N USB_HDMI_WiFi_BT_Ethernet_LCD_HTX2P R
  XR43 USB_HDMI_WiFi_BT_Ethernet_LCD_HTX1P USB_HDMI_WiFi_BT_Ethernet_LCD_HTX1N R
  XR44 USB_HDMI_WiFi_BT_Ethernet_LCD_HTX0N USB_HDMI_WiFi_BT_Ethernet_LCD_HTX0P R
  XR45 USB_HDMI_WiFi_BT_Ethernet_LCD_HTXCP USB_HDMI_WiFi_BT_Ethernet_LCD_HTXCN R
  XC79 GND _3.3VD C
  XUSB_OTG1 GND GND GND GND _5V_USBOTG USB0_D_N USB0_D_P USB_HDMI_WiFi_BT_Ethernet_LCD_USB0_ID GND USB-MINI
  XR37 USB_HDMI_WiFi_BT_Ethernet_LCD_USB0_ID _3.3V R
  XU6 Net__C68_Pad2_ GND Net__R41_Pad2_ USB0_DRV _5V SY6280AAC(SOT23-5)
  XL6 Net__C68_Pad2_ _5V_USBOTG L
  XC67 _5V_USBOTG GND C
  XC70 GND Net__C68_Pad2_ C
  XC69 GND Net__C68_Pad2_ C
  XC68 GND Net__C68_Pad2_ C
  XR41 GND Net__R41_Pad2_ R
  XR38 USB_HDMI_WiFi_BT_Ethernet_LCD_USB0_VBUSDET Net__C68_Pad2_ R
  XR42 GND USB_HDMI_WiFi_BT_Ethernet_LCD_USB0_VBUSDET R
  XC72 GND USB_HDMI_WiFi_BT_Ethernet_LCD_USB0_VBUSDET C
  XR40 GND USB0_DRV R
  XC71 _5V GND C
  XU9 Net__C75_Pad2_ GND Net__R49_Pad2_ USB1_DRV _5V SY6280AAC(SOT23-5)
  XL8 Net__C75_Pad2_ Net__C74_Pad1_ L
  XC74 Net__C74_Pad1_ GND C
  XC77 GND Net__C75_Pad2_ C
  XC76 GND Net__C75_Pad2_ C
  XC75 GND Net__C75_Pad2_ C
  XR49 GND Net__R49_Pad2_ R
  XR48 GND USB1_DRV R
  XC78 _5V GND C
  XC73 GND _3.3V C
  XC110 GND _3.3VWiFiIO C
  XU11 GND Net__U11_Pad10_ Net__U11_Pad11_ USB_HDMI_WiFi_BT_Ethernet_LCD_WL_PMU_EN USB_HDMI_WiFi_BT_Ethernet_LCD_WL_WAKE_AP USB_HDMI_WiFi_BT_Ethernet_LCD_WL_SDIO_D2 USB_HDMI_WiFi_BT_Ethernet_LCD_WL_SDIO_D3 USB_HDMI_WiFi_BT_Ethernet_LCD_WL_SDIO_CMD Net__R54_Pad1_ USB_HDMI_WiFi_BT_Ethernet_LCD_WL_SDIO_D0 USB_HDMI_WiFi_BT_Ethernet_LCD_WL_SDIO_D1 Net__C105_Pad1_ GND Net__U11_Pad21_ _3.3VWiFiIO Net__U11_Pad23_ Net__R60_Pad1_ USB_HDMI_WiFi_BT_Ethernet_LCD_BT_PCM_DOUT USB_HDMI_WiFi_BT_Ethernet_LCD_BT_PCM_CLK USB_HDMI_WiFi_BT_Ethernet_LCD_BT_PCM_DIN USB_HDMI_WiFi_BT_Ethernet_LCD_BT_PCM_SYNC Net__U11_Pad29_ Net__U11_Pad3_ Net__U11_Pad30_ GND Net__U11_Pad32_ GND USB_HDMI_WiFi_BT_Ethernet_LCD_BT_RST_N Net__U11_Pad35_ GND Net__U11_Pad37_ Net__U11_Pad38_ Net__U11_Pad39_ Net__U11_Pad4_ Net__U11_Pad40_ GND USB_HDMI_WiFi_BT_Ethernet_LCD_BT_UART_TX USB_HDMI_WiFi_BT_Ethernet_LCD_BT_UART_RX USB_HDMI_WiFi_BT_Ethernet_LCD_BT_UART_CTS Net__U11_Pad5_ USB_HDMI_WiFi_BT_Ethernet_LCD_AP_WAKE_BT USB_HDMI_WiFi_BT_Ethernet_LCD_BT_WAKE_AP Net__U11_Pad8_ _3.3V RTL8723BS(ComboModule)
  XR54 Net__R54_Pad1_ USB_HDMI_WiFi_BT_Ethernet_LCD_WL_SDIO_CLK R
  XRM9 _3.3VWiFiIO USB_HDMI_WiFi_BT_Ethernet_LCD_WL_SDIO_D0 _3.3VWiFiIO USB_HDMI_WiFi_BT_Ethernet_LCD_WL_SDIO_D3 _3.3VWiFiIO USB_HDMI_WiFi_BT_Ethernet_LCD_WL_SDIO_D2 _3.3VWiFiIO USB_HDMI_WiFi_BT_Ethernet_LCD_WL_PMU_EN RA1206_(4x0603)_4B8_Smashed
  XC92 GND _3.3VWiFiIO C
  XC91 GND _3.3VWiFiIO C
  XC90 GND _3.3V C
  XC89 GND _3.3V C
  XC109 VCC_PL GND C
  XC105 Net__C105_Pad1_ Net__C105_Pad2_ C
  XC106 GND Net__C105_Pad2_ C
  XC107 GND Net__C107_Pad2_ C
  XANT1 Net__ANT1_Pad1_ GND WIFI_ANT_ESP8266
  XRM12 _3.3VWiFiIO USB_HDMI_WiFi_BT_Ethernet_LCD_WL_SDIO_CMD _3.3VWiFiIO USB_HDMI_WiFi_BT_Ethernet_LCD_BT_RST_N _3.3VWiFiIO USB_HDMI_WiFi_BT_Ethernet_LCD_WL_SDIO_D1 _3.3VWiFiIO USB_HDMI_WiFi_BT_Ethernet_LCD_BT_UART_RX RA1206_(4x0603)_4B8_Smashed
  XR61 AP_CK32KO _3.3VWiFiIO R
  XC80 _3.3V GND C
  XR70 TWI0_SCK _3.3V R
  XR71 TWI0_SDA _3.3V R
  XLCD_CON1 GND _5V USB_HDMI_WiFi_BT_Ethernet_LCD_GTXD3_LCD_D21 USB_HDMI_WiFi_BT_Ethernet_LCD_GTXD2_LCD_D22 USB_HDMI_WiFi_BT_Ethernet_LCD_GTXD1_LCD_D23 GND GND USB_HDMI_WiFi_BT_Ethernet_LCD_LCD_D10 USB_HDMI_WiFi_BT_Ethernet_LCD_LCD_D11 USB_HDMI_WiFi_BT_Ethernet_LCD_GRXD3_LCD_D12 USB_HDMI_WiFi_BT_Ethernet_LCD_GRXD2_LCD_D13 USB_HDMI_WiFi_BT_Ethernet_LCD_GRXD1_LCD_D14 GND USB_HDMI_WiFi_BT_Ethernet_LCD_GRXD0_LCD_D15 GND GND USB_HDMI_WiFi_BT_Ethernet_LCD_LCD_D2 USB_HDMI_WiFi_BT_Ethernet_LCD_LCD_D3 USB_HDMI_WiFi_BT_Ethernet_LCD_LCD_D4 USB_HDMI_WiFi_BT_Ethernet_LCD_LCD_D5 USB_HDMI_WiFi_BT_Ethernet_LCD_LCD_D6 USB_HDMI_WiFi_BT_Ethernet_LCD_LCD_D7 USB_HDMI_WiFi_BT_Ethernet_LCD_GTXCTL_LCD_HSYNC _3.3V USB_HDMI_WiFi_BT_Ethernet_LCD_GCLKIN_LCD_VSYNC USB_HDMI_WiFi_BT_Ethernet_LCD_GTXD0_LCD_CLK USB_HDMI_WiFi_BT_Ethernet_LCD_GTXCK_LCD_DE PH10 PH11 USB_HDMI_WiFi_BT_Ethernet_LCD_GMDIO_LCD_PWR USB_HDMI_WiFi_BT_Ethernet_LCD_GMDC_LCD_PWM USB_HDMI_WiFi_BT_Ethernet_LCD_PH7_CTP_INT USB_HDMI_WiFi_BT_Ethernet_LCD_PH8_CTP_RST TWI0_SCK GND TWI0_SDA GND GND USB_HDMI_WiFi_BT_Ethernet_LCD_GRXCK_LCD_D18 USB_HDMI_WiFi_BT_Ethernet_LCD_GRXCTL_LCD_D19 USB_HDMI_WiFi_BT_Ethernet_LCD_LCD_D20 LCD-ML40YA-V36P-2X20-LF
  XR99 _3.3V USB1_DRV R
  XUSB1 GND GND Net__C74_Pad1_ USB_HDMI_WiFi_BT_Ethernet_LCD_USB1_DM USB_HDMI_WiFi_BT_Ethernet_LCD_USB1_DP GND USB_A_VERTICAL
  XU15 USB_HDMI_WiFi_BT_Ethernet_LCD_VDD33 USB_HDMI_WiFi_BT_Ethernet_LCD_MDI_3___0 USB_HDMI_WiFi_BT_Ethernet_LCD_MDI_3__ USB_HDMI_WiFi_BT_Ethernet_LCD_VDD33 Net__U15_Pad13_ Net__C204_Pad2_ Net__R113_Pad2_ USB_HDMI_WiFi_BT_Ethernet_LCD_VDD33 Net__R111_Pad2_ Net__C204_Pad2_ USB_HDMI_WiFi_BT_Ethernet_LCD_GTXD0_LCD_CLK USB_HDMI_WiFi_BT_Ethernet_LCD_MDI_0___0 USB_HDMI_WiFi_BT_Ethernet_LCD_GTXD1_LCD_D23 USB_HDMI_WiFi_BT_Ethernet_LCD_GTXD2_LCD_D22 USB_HDMI_WiFi_BT_Ethernet_LCD_GTXD3_LCD_D21 Net__C204_Pad2_ USB_HDMI_WiFi_BT_Ethernet_LCD_GTXCK_LCD_DE USB_HDMI_WiFi_BT_Ethernet_LCD_GTXCTL_LCD_HSYNC Net__C204_Pad2_ Net__RM15_Pad4.1_ Net__RM15_Pad3.1_ GND USB_HDMI_WiFi_BT_Ethernet_LCD_MDI_0__ Net__C204_Pad2_ Net__RM15_Pad2.1_ Net__RM15_Pad1.1_ Net__R105_Pad2_ USB_HDMI_WiFi_BT_Ethernet_LCD_VDD33 Net__R107_Pad1_ USB_HDMI_WiFi_BT_Ethernet_LCD_GMDC_LCD_PWM USB_HDMI_WiFi_BT_Ethernet_LCD_GMDIO_LCD_PWR Net__R119_Pad1_ Net__C204_Pad2_ Net__C207_Pad2_ USB_HDMI_WiFi_BT_Ethernet_LCD_VDD33 Net__R109_Pad2_ Net__C211_Pad2_ Net__U15_Pad43_ Net__C207_Pad2_ Net__C213_Pad2_ Net__C212_Pad2_ Net__U15_Pad47_ Net__R115_Pad1_ GND USB_HDMI_WiFi_BT_Ethernet_LCD_MDI_1__ USB_HDMI_WiFi_BT_Ethernet_LCD_MDI_1___0 USB_HDMI_WiFi_BT_Ethernet_LCD_MDI_2__ USB_HDMI_WiFi_BT_Ethernet_LCD_MDI_2___0 Net__C207_Pad2_ KSZ9031RNXCC(QFN48_1DRILL(PADPITCH-0.5MM))
  XRM8 USB_HDMI_WiFi_BT_Ethernet_LCD_VDD33 Net__RM15_Pad1.1_ USB_HDMI_WiFi_BT_Ethernet_LCD_VDD33 Net__RM15_Pad2.1_ USB_HDMI_WiFi_BT_Ethernet_LCD_VDD33 Net__RM15_Pad3.1_ USB_HDMI_WiFi_BT_Ethernet_LCD_VDD33 Net__RM15_Pad4.1_ RA1206_(4x0603)_4B8_Smashed
  XR105 USB_HDMI_WiFi_BT_Ethernet_LCD_GRXCTL_LCD_D19 Net__R105_Pad2_ R
  XR106 USB_HDMI_WiFi_BT_Ethernet_LCD_VDD33 Net__R105_Pad2_ R
  XR107 Net__R107_Pad1_ GND R
  XC198 USB_HDMI_WiFi_BT_Ethernet_LCD_GRXCK_LCD_D18 Net__C198_Pad2_ C
  XR108 USB_HDMI_WiFi_BT_Ethernet_LCD_GMDIO_LCD_PWR USB_HDMI_WiFi_BT_Ethernet_LCD_VDD33 R
  XR109 USB_HDMI_WiFi_BT_Ethernet_LCD_GCLKIN_LCD_VSYNC Net__R109_Pad2_ R
  XR110 USB_HDMI_WiFi_BT_Ethernet_LCD_VDD33 Net__R109_Pad2_ R
  XR111 USB_HDMI_WiFi_BT_Ethernet_LCD_VDD33 Net__R111_Pad2_ R
  XR112 USB_HDMI_WiFi_BT_Ethernet_LCD_PHYAD0 Net__R111_Pad2_ R
  XR113 USB_HDMI_WiFi_BT_Ethernet_LCD_PHYAD1 Net__R113_Pad2_ R
  XR114 GND Net__R113_Pad2_ R
  XLAN1 USB_HDMI_WiFi_BT_Ethernet_LCD_MDI_0___0 USB_HDMI_WiFi_BT_Ethernet_LCD_MDI_3__ USB_HDMI_WiFi_BT_Ethernet_LCD_VDD33 USB_HDMI_WiFi_BT_Ethernet_LCD_PHYAD1 USB_HDMI_WiFi_BT_Ethernet_LCD_VDD33 USB_HDMI_WiFi_BT_Ethernet_LCD_PHYAD0 USB_HDMI_WiFi_BT_Ethernet_LCD_MDI_0__ USB_HDMI_WiFi_BT_Ethernet_LCD_MDI_1__ USB_HDMI_WiFi_BT_Ethernet_LCD_MDI_1___0 Net__C199_Pad2_ Net__C200_Pad2_ USB_HDMI_WiFi_BT_Ethernet_LCD_MDI_2__ USB_HDMI_WiFi_BT_Ethernet_LCD_MDI_2___0 USB_HDMI_WiFi_BT_Ethernet_LCD_MDI_3___0 Net__C196_Pad2_ Net__C196_Pad2_ TM211Q01FM22
  XC199 GND Net__C199_Pad2_ C
  XC200 GND Net__C200_Pad2_ C
  XC196 GND Net__C196_Pad2_ C
  XL21 USB_HDMI_WiFi_BT_Ethernet_LCD_VDD33 _3.3V L
  XC201 USB_HDMI_WiFi_BT_Ethernet_LCD_VDD33 GND C
  XC216 GND USB_HDMI_WiFi_BT_Ethernet_LCD_VDD33 C
  XC214 GND Net__C207_Pad2_ C
  XC207 GND Net__C207_Pad2_ C
  XC215 GND Net__C207_Pad2_ C
  XC202 USB_HDMI_WiFi_BT_Ethernet_LCD_VDD33 GND C
  XC217 GND USB_HDMI_WiFi_BT_Ethernet_LCD_VDD33 C
  XC203 GND USB_HDMI_WiFi_BT_Ethernet_LCD_VDD33 C
  XC204 GND Net__C204_Pad2_ C
  XC208 GND Net__C204_Pad2_ C
  XC205 GND Net__C204_Pad2_ C
  XC209 GND Net__C204_Pad2_ C
  XC206 GND Net__C204_Pad2_ C
  XC210 GND Net__C204_Pad2_ C
  XR115 Net__R115_Pad1_ GND R
  XR116 Net__C211_Pad2_ USB_HDMI_WiFi_BT_Ethernet_LCD_VDD33 R
  XR117 Net__C211_Pad2_ USB_HDMI_WiFi_BT_Ethernet_LCD_EPHY_RST_ R
  XR118 Net__C211_Pad2_ AP_RESET_ R
  XR119 Net__R119_Pad1_ USB_HDMI_WiFi_BT_Ethernet_LCD_VDD33 R
  XC211 GND Net__C211_Pad2_ C
  XC212 GND Net__C212_Pad2_ C
  XC213 GND Net__C213_Pad2_ C
  XL23 Net__C207_Pad2_ USB_HDMI_WiFi_BT_Ethernet_LCD_1.25_EXT L
  XL24 Net__C204_Pad2_ USB_HDMI_WiFi_BT_Ethernet_LCD_1.25_EXT L
  XC218 Net__C218_Pad1_ GND C
  XVR1 GND USB_HDMI_WiFi_BT_Ethernet_LCD_1.25_EXT Net__C218_Pad1_ AMS1117-ADJ
  XR120 USB_HDMI_WiFi_BT_Ethernet_LCD_1.25_EXT GND R
  XC219 USB_HDMI_WiFi_BT_Ethernet_LCD_1.25_EXT GND C
  XPHYRST1 GND Net__C211_Pad2_ JP1E
  XD5 Net__C218_Pad1_ _3.3V D
  X_1.25_EXT1 USB_HDMI_WiFi_BT_Ethernet_LCD_1.25_EXT TESTPAD
  XRM15 Net__RM15_Pad1.1_ USB_HDMI_WiFi_BT_Ethernet_LCD_GRXD0_LCD_D15 Net__RM15_Pad2.1_ USB_HDMI_WiFi_BT_Ethernet_LCD_GRXD1_LCD_D14 Net__RM15_Pad3.1_ USB_HDMI_WiFi_BT_Ethernet_LCD_GRXD2_LCD_D13 Net__RM15_Pad4.1_ USB_HDMI_WiFi_BT_Ethernet_LCD_GRXD3_LCD_D12 RA1206_(4x0603)_4B8_Smashed
  XRM1 USB_HDMI_WiFi_BT_Ethernet_LCD_GTXD1_LCD_D23 Net__RM1_Pad1.2_ USB_HDMI_WiFi_BT_Ethernet_LCD_GTXD0_LCD_CLK Net__RM1_Pad2.2_ USB_HDMI_WiFi_BT_Ethernet_LCD_GTXD2_LCD_D22 Net__RM1_Pad3.2_ USB_HDMI_WiFi_BT_Ethernet_LCD_GTXD3_LCD_D21 Net__RM1_Pad4.2_ RA1206_(4x0603)_4B8_Smashed
  XR72 Net__R72_Pad1_ USB_HDMI_WiFi_BT_Ethernet_LCD_GTXCTL_LCD_HSYNC R
  XL9 Net__C88_Pad2_ USB_HDMI_WiFi_BT_Ethernet_LCD_GTXCK_LCD_DE L
  XL7 Net__C198_Pad2_ GND L
  XC93 GND USB_HDMI_WiFi_BT_Ethernet_LCD_GCLKIN_LCD_VSYNC C
  XL10 Net__C107_Pad2_ Net__C105_Pad2_ L
  XC88 GND Net__C88_Pad2_ C
  XU4 _3.3V _3.3V _3.3V GND TWI1_SDA TWI1_SCK GND _3.3V AT24C16BN-SH(SO-8_150mil)
  XC39 _3.3V GND C
  XANT2 Net__ANT2_Pad1_ GND WIFI_ANT_ESP8266
  XR60 Net__R60_Pad1_ AP_CK32KO R
  XR17 Net__ANT2_Pad1_ Net__C107_Pad2_ R
  XR16 Net__ANT1_Pad1_ Net__C107_Pad2_ R
  XR18 USB_HDMI_WiFi_BT_Ethernet_LCD_GRXCK_LCD_D18 Net__R107_Pad1_ R
  XR19 Net__R19_Pad1_ USB_HDMI_WiFi_BT_Ethernet_LCD_GTXCK_LCD_DE R
  XQ4 Net__C212_Pad2_ Net__C213_Pad2_ GND Crystal_GND
  XD3 Net__D3_Pad1_ _5V D_Schottky
  XTVS1 USB_HDMI_WiFi_BT_Ethernet_LCD_MDI_0___0 USB_HDMI_WiFi_BT_Ethernet_LCD_MDI_0___0 GND USB_HDMI_WiFi_BT_Ethernet_LCD_MDI_1__ USB_HDMI_WiFi_BT_Ethernet_LCD_MDI_1___0 USB_HDMI_WiFi_BT_Ethernet_LCD_MDI_0__ ESDS314DBVR(SOT-23-5)
  XTVS2 USB_HDMI_WiFi_BT_Ethernet_LCD_MDI_2___0 USB_HDMI_WiFi_BT_Ethernet_LCD_MDI_2___0 GND USB_HDMI_WiFi_BT_Ethernet_LCD_MDI_3__ USB_HDMI_WiFi_BT_Ethernet_LCD_MDI_3___0 USB_HDMI_WiFi_BT_Ethernet_LCD_MDI_2__ ESDS314DBVR(SOT-23-5)
  XU14 Power_Supply__Extensions_and_MiPi_DSI_1.8V_DVDD_CSI Net__L20_Pad1_ IPS GND _3.3VWiFiIO Power_Supply__Extensions_and_MiPi_DSI_2.8V_AVDD_CSI IPS Power_Supply__Extensions_and_MiPi_DSI_3.3V_MIPI _3.3VD Net__C125_Pad2_ IPS Net__C174_Pad2_ _3.3V Net__L14_Pad1_ IPS Net__U14_Pad23_ Net__U14_Pad24_ GND Net__R86_Pad1_ Net__R87_Pad1_ VCC_PE VCC_PL _1.2V_HSIC Net__R83_Pad1_ _3.0VA IPS Net__C182_Pad2_ Net__C151_Pad1_ Net__C149_Pad1_ Net__L17_Pad1_ Net__L17_Pad1_ IPS IPS IPS IPS VDDFB_CPUX VDDFB_CPUX Net__L15_Pad1_ Net__L15_Pad1_ GND AP_RESET_ PMU_SCK PMU_SDA _3.0V_RTC _1.1V_CPUS Net__C181_Pad2_ USB0_DRV Net__T1_Pad3_ Net__R82_Pad1_ _5V_USBOTG IPS IPS _5V_EXT _5V_EXT GND IPS Net__C177_Pad2_ AP_NMI_ Power_Supply__Extensions_and_MiPi_DSI_DC5SET Net__C135_Pad1_ VBAT Net__L18_Pad2_ IPS IPS _1.8V GND Net__L19_Pad1_ _1.5V _1.1V_SYS AXP803
  XC177 GND Net__C177_Pad2_ C
  XR91 Net__PWRON1_Pad1_ Net__C177_Pad2_ R
  XC121 _5V_EXT GND C
  XPWR1 _5V_EXT GND GND PWR-JAKPWR_JACK_UNI_MILLING
  XFUSE2 _5V_EXT _5V_EXT FSMD035
  XC118 GND _5V_EXT C
  XC119 GND _5V_EXT C
  XC124 _5V_USBOTG GND C
  XC128 IPS GND C
  XL14 Net__L14_Pad1_ _3.3V L
  XC122 GND _3.3V C
  XC125 GND Net__C125_Pad2_ C
  XC126 GND IPS C
  XL15 Net__L15_Pad1_ _1.1V_CPUX L
  XC129 GND _1.1V_CPUX C
  XC131 GND _1.1V_CPUX C
  XC133 GND IPS C
  XL17 Net__L17_Pad1_ _1.1V_CPUX L
  XC136 GND _1.1V_CPUX C
  XC139 GND _1.1V_CPUX C
  XC145 GND IPS C
  XL19 Net__L19_Pad1_ _1.5V L
  XC150 GND _1.5V C
  XC153 GND IPS C
  XR84 GND Power_Supply__Extensions_and_MiPi_DSI_DC5SET R
  XL20 Net__L20_Pad1_ _1.1V_SYS L
  XC154 GND _1.1V_SYS C
  XC157 GND IPS C
  XC159 GND IPS C
  XC161 GND _3.3VD C
  XC162 GND Power_Supply__Extensions_and_MiPi_DSI_3.3V_MIPI C
  XC164 GND Power_Supply__Extensions_and_MiPi_DSI_2.8V_AVDD_CSI C
  XC165 GND _3.3VWiFiIO C
  XC167 GND IPS C
  XC176 GND IPS C
  XC169 IPS GND C
  XT1 Net__C135_Pad1_ Net__C135_Pad1_ Net__T1_Pad3_ IPS Net__C135_Pad1_ Net__C135_Pad1_ Net__C135_Pad1_ IPS WPM1481
  XR78 Net__C135_Pad1_ VBAT R
  XC135 Net__C135_Pad1_ VBAT C
  XL18 Net__C135_Pad1_ Net__L18_Pad2_ L
  XC144 Net__C135_Pad1_ GND C
  XC138 Net__C135_Pad1_ GND C
  XC147 IPS GND C
  XCHGLED1 Net__CHGLED1_Pad1_ IPS LED
  XR82 Net__R82_Pad1_ Net__CHGLED1_Pad1_ R
  XR83 Net__R83_Pad1_ GND R
  XC149 Net__C149_Pad1_ GND C
  XC151 Net__C151_Pad1_ GND C
  XC152 _3.0V_RTC GND C
  XR85 AP_NMI_ _3.0V_RTC R
  XR86 Net__R86_Pad1_ USB0_D_P R
  XR87 Net__R87_Pad1_ USB0_D_N R
  XR88 PMU_SCK VCC_PL R
  XR90 PMU_SDA VCC_PL R
  XC173 VCC_PL GND C
  XC175 _3.0VA GND C
  XC171 VCC_PE GND C
  XPWRON1 Net__PWRON1_Pad1_ GND T1107A(6x3,8x2,5MM)
  XC156 GND AP_RESET_ C
  XR89 Net__R89_Pad1_ AP_RESET_ R
  XRESET1 Net__R89_Pad1_ GND T1107A(6x3,8x2,5MM)
  XC160 GND _1.1V_SYS C
  XC163 GND _1.1V_SYS C
  XC155 GND _1.1V_SYS C
  XC158 GND _1.1V_SYS C
  XC166 GND _1.1V_SYS C
  XC168 GND _1.1V_SYS C
  XC142 GND _1.1V_CPUX C
  XC137 GND _1.1V_CPUX C
  XC123 GND _1.1V_CPUX C
  XC148 GND _1.1V_CPUX C
  XC146 GND _1.1V_CPUX C
  XC127 GND _1.1V_CPUX C
  XC130 GND _1.1V_CPUX C
  XC132 GND _1.1V_CPUX C
  XC134 GND _1.1V_CPUX C
  XC117 GND _1.1V_CPUS C
  XC120 GND _1.1V_CPUS C
  XC179 GND _1.1V_CPUS C
  XC115 GND _3.3V C
  XC116 GND _3.3V C
  XC185 Net__C185_Pad1_ GND C
  XC187 Net__C187_Pad1_ GND C
  XR94 Net__R94_Pad1_ Net__C185_Pad1_ R
  XQ2 Net__C183_Pad1_ Net__C184_Pad1_ Crystal
  XC183 Net__C183_Pad1_ GND C
  XC184 Net__C184_Pad1_ GND C
  XR93 Net__C183_Pad1_ Net__C184_Pad1_ R
  XR96 Net__R96_Pad1_ GND R
  XR97 Net__R97_Pad1_ GND R
  XR98 Net__R98_Pad1_ GND R
  XC193 GND KEYADC C
  XUBOOT1 UBOOT GND T1107A(6x3,8x2,5MM)
  XC178 GND _1.2V_HSIC C
  XC186 GND _3.3V C
  XC188 GND Net__C188_Pad2_ C
  XC190 GND _3.0V_RTC C
  XC189 GND _3.0V_RTC C
  XC191 GND _3.0VA C
  XC192 GND Net__C192_Pad2_ C
  XDBG_UART1 Net__DBG_UART1_Pad1_ Net__D4_Pad1_ GND CON3
  XD4 Net__D4_Pad1_ Net__D4_Pad2_ D_Schottky
  XR95 Net__D4_Pad2_ _3.3V R
  XC170 GND _1.8V C
  XUEXT1 _3.3V Power_Supply__Extensions_and_MiPi_DSI_UEXT_CS GND UART3_TX UART3_RX TWI1_SCK TWI1_SDA Power_Supply__Extensions_and_MiPi_DSI_UEXT_MISO Power_Supply__Extensions_and_MiPi_DSI_UEXT_MOSI Power_Supply__Extensions_and_MiPi_DSI_UEXT_CLK BH10S
  XR75 _3.3V TWI1_SCK R
  XR76 _3.3V UART3_RX R
  XR77 _3.3V TWI1_SDA R
  XD1 _5V_EXT GND SMBJ6.0A
  XPWRLED1 GND Net__PWRLED1_Pad2_ LED
  XR74 _5V_EXT Net__PWRLED1_Pad2_ R
  X_5V_E1 _5V_EXT _5V SJ
  XC172 GND Power_Supply__Extensions_and_MiPi_DSI_1.8V_DVDD_CSI C
  XC174 GND Net__C174_Pad2_ C
  XC181 GND Net__C181_Pad2_ C
  XC182 GND Net__C182_Pad2_ C
  XR92 Power_Supply__Extensions_and_MiPi_DSI_DC5SET Net__C181_Pad2_ R
  XLIPO_BAT1 VBAT GND CON2
  XC180 GND VBAT C
  XGPIO1 _5V Power_Supply__Extensions_and_MiPi_DSI_PB0 Power_Supply__Extensions_and_MiPi_DSI_PE3 Power_Supply__Extensions_and_MiPi_DSI_PB1 Power_Supply__Extensions_and_MiPi_DSI_PE4 Power_Supply__Extensions_and_MiPi_DSI_PB2 Power_Supply__Extensions_and_MiPi_DSI_PE5 Power_Supply__Extensions_and_MiPi_DSI_PB3 Power_Supply__Extensions_and_MiPi_DSI_PE6 Power_Supply__Extensions_and_MiPi_DSI_PB4 Power_Supply__Extensions_and_MiPi_DSI_PE7 GND PC4 Power_Supply__Extensions_and_MiPi_DSI_PE8 PC7 Power_Supply__Extensions_and_MiPi_DSI_PE9 PL7 Power_Supply__Extensions_and_MiPi_DSI_PE10 PL8 Power_Supply__Extensions_and_MiPi_DSI_PE11 PL9 Power_Supply__Extensions_and_MiPi_DSI_PE12 _3.3V PL10 Power_Supply__Extensions_and_MiPi_DSI_PE13 PL11 Power_Supply__Extensions_and_MiPi_DSI_PE14 PL12 Power_Supply__Extensions_and_MiPi_DSI_PE15 Power_Supply__Extensions_and_MiPi_DSI_1.8V_DVDD_CSI Power_Supply__Extensions_and_MiPi_DSI_PE16__POWERON Power_Supply__Extensions_and_MiPi_DSI_2.8V_AVDD_CSI Power_Supply__Extensions_and_MiPi_DSI_PE17__GPIO_LED AP_RESET_ VCC_PE Power_Supply__Extensions_and_MiPi_DSI_PE0 UBOOT Power_Supply__Extensions_and_MiPi_DSI_PE1 KEYADC Power_Supply__Extensions_and_MiPi_DSI_PE2 ML40YA-V36P-2X20-LF
  XMIPI_DSI1 GND GND TWI0_SCK TWI0_SDA GND Power_Supply__Extensions_and_MiPi_DSI_3.3V_MIPI Power_Supply__Extensions_and_MiPi_DSI_3.3V_MIPI Net__MIPI_DSI1_Pad16_ Net__MIPI_DSI1_Pad17_ GND Net__MIPI_DSI1_Pad19_ Power_Supply__Extensions_and_MiPi_DSI_DSI_D1N Net__MIPI_DSI1_Pad20_ Power_Supply__Extensions_and_MiPi_DSI_DSI_D1P GND Power_Supply__Extensions_and_MiPi_DSI_DSI_CKN Power_Supply__Extensions_and_MiPi_DSI_DSI_CKP GND Power_Supply__Extensions_and_MiPi_DSI_DSI_D0N Power_Supply__Extensions_and_MiPi_DSI_DSI_D0P GPH127SMT-02X10(PA-V16X-2X10-LF)
  XC195 GND _3.3V C
  XC194 GND Net__3.3V_VCC_PE_2.8V1_Pad2_ C
  X_3.3V_VCC_PE_2.8V1 VCC_PE Net__3.3V_VCC_PE_2.8V1_Pad2_ _3.3V SJ2W_Closed(1-2)
  XR79 _3.3V Power_Supply__Extensions_and_MiPi_DSI_UEXT_CS R
  XR102 Power_Supply__Extensions_and_MiPi_DSI_PE15 Net__3.3V_VCC_PE_2.8V1_Pad2_ R
  XR101 Power_Supply__Extensions_and_MiPi_DSI_PE14 Net__3.3V_VCC_PE_2.8V1_Pad2_ R
  XHSIC1 Net__HSIC1_Pad1_ Net__HSIC1_Pad2_ Net__HSIC1_Pad3_ GND CON4
  XHSIC_E1 _1.2V_HSIC Net__HSIC1_Pad1_ SJ
  XC197 _1.2V_HSIC GND C
  XR103 _3.0VA KEYADC R
  XR104 _3.0V_RTC AP_RESET_ R
  XGPIO_LED1 GND Net__GPIO_LED1_Pad2_ LED
  XR58 Power_Supply__Extensions_and_MiPi_DSI_PE17__GPIO_LED Net__GPIO_LED1_Pad2_ R
  X_3.3V1 _3.3V TESTPAD
  X_1.1V_CPUX1 _1.1V_CPUX TESTPAD
  XDDR_VCC1 _1.5V TESTPAD
  X_1.1V_SYS1 _1.1V_SYS TESTPAD
  X_3.3VD1 _3.3VD TESTPAD
  X_3.3VWiFiIO1 _3.3VWiFiIO TESTPAD
  X_3.3V_MIPI1 Power_Supply__Extensions_and_MiPi_DSI_3.3V_MIPI TESTPAD
  X_5V_USBOTG1 _5V_USBOTG TESTPAD
  XIPS1 IPS TESTPAD
  X_3.0V_RTC1 _3.0V_RTC TESTPAD
  XVCC_PC1 VCC_PC TESTPAD
  X_1.8V1 _1.8V TESTPAD
  X_1.1V_CPUS1 _1.1V_CPUS TESTPAD
  X_3.0VA1 _3.0VA TESTPAD
  XVCC_PL1 VCC_PL TESTPAD
  XGND1 GND TESTPAD
  XR65 Power_Supply__Extensions_and_MiPi_DSI_PE16__POWERON Power_Supply__Extensions_and_MiPi_DSI_PE16 R
  XR28 Power_Supply__Extensions_and_MiPi_DSI_PE16__POWERON Net__C177_Pad2_ R
  XPWR_PC1 _3.3V VCC_PC _1.8V SJ2W
  XR121 Power_Supply__Extensions_and_MiPi_DSI_UEXT_MISO SPI0_MISO R
  XR122 Power_Supply__Extensions_and_MiPi_DSI_UEXT_CLK SPI0_CLK R
  XR123 SPI0_MOSI Power_Supply__Extensions_and_MiPi_DSI_UEXT_MOSI R
  XR124 SPI0_CS Power_Supply__Extensions_and_MiPi_DSI_UEXT_CS R
  XR73 PH10 Power_Supply__Extensions_and_MiPi_DSI_UEXT_CS R
  XR125 Net__MIPI_DSI1_Pad17_ Power_Supply__Extensions_and_MiPi_DSI_DSI_D3P R
  XR126 Net__MIPI_DSI1_Pad19_ Power_Supply__Extensions_and_MiPi_DSI_DSI_D2N R
  XR130 Power_Supply__Extensions_and_MiPi_DSI_DSI_D2P Net__MIPI_DSI1_Pad20_ R
  XR129 Power_Supply__Extensions_and_MiPi_DSI_DSI_D3N Net__MIPI_DSI1_Pad16_ R
  XR128 Net__MIPI_DSI1_Pad19_ Power_Supply__Extensions_and_MiPi_DSI_MIPI_DSI_EN R
  XR127 Net__MIPI_DSI1_Pad17_ Power_Supply__Extensions_and_MiPi_DSI_MIPI_DSI_RST R
  XR132 Power_Supply__Extensions_and_MiPi_DSI_MIPI_DSI_BKL Net__MIPI_DSI1_Pad20_ R
  XR131 IPS Net__MIPI_DSI1_Pad16_ R
  XQ3 Net__C185_Pad1_ Net__C187_Pad1_ GND Crystal_GND
  XU16 Net__FET3_Pad1_ GND _5V_EXT VDA2710NTA(SOT-23)
  XFET4 Net__FET3_Pad1_ GND Net__FET2_Pad1_ N-MOS+DIOD_Small
  XR20 Net__FET3_Pad1_ _5V_EXT R
  XR24 _5V Net__FET2_Pad1_ R
  XFET2 Net__FET2_Pad1_ _5V _5V_EXT P-MOS+DIOD
  XR22 GND Net__FET3_Pad1_ R
  XFET3 Net__FET3_Pad1_ _5V Net__C143_Pad2_ P-MOS+DIOD
  XC143 GND Net__C143_Pad2_ C
  XC140 GND IPS C
  XR81 Net__R80_Pad2_ GND R
  XR80 Net__C143_Pad2_ Net__R80_Pad2_ R
  XD2 Net__C143_Pad2_ Net__D2_Pad2_ D_Schottky
  XL16 IPS Net__D2_Pad2_ L
  XC141 GND IPS C
  XU13 Net__D2_Pad2_ GND Net__R80_Pad2_ _3.3V IPS Net__U13_Pad6_ MT3608(SOT23-6)
.ends A64-OlinuXino_Rev_H

*--- Subcircuit Definitions ---
.subckt C 1 2
* Stub for C
.ends

.subckt R 1 2
* Stub for R
.ends

.subckt H5TQ2G63BFR_MEM4G16D3EABG-125--H5TC8G63AMR-PBA_K4B8G1646Q-MYK0(FBGA-96_512MX16_DDR3-1600_11-11-11) A1 A2 A3 A7 A8 A9 B1 B2 B3 B7 B8 B9 C1 C2 C3 C7 C8 C9 D1 D2 D3 D7 D8 D9 E1 E2 E3 E7 E8 E9 F1 F2 F3 F7 F8 F9 G1 G2 G3 G7 G8 G9 H1 H2 H3 H7 H8 H9 J1 J2 J3 J7 J8 J9 K1 K2 K3 K7 K8 K9 L1 L2 L3 L7 L8 L9 M1 M2 M3 M7 M8 M9 N1 N2 N3 N7 N8 N9 P1 P2 P3 P7 P8 P9 R1 R2 R3 R7 R8 R9 T1 T2 T3 T7 T8 T9
* Stub for H5TQ2G63BFR_MEM4G16D3EABG-125--H5TC8G63AMR-PBA_K4B8G1646Q-MYK0(FBGA-96_512MX16_DDR3-1600_11-11-11)
.ends

.subckt AllWinner-A64(FBGA396) A1 A11 A13 A14 A16 A17 A19 A2 A20 A22 A23 A4 A5 A7 A8 AA1 AA10 AA11 AA12 AA13 AA14 AA15 AA16 AA17 AA18 AA19 AA20 AA21 AA22 AA3 AA5 AA6 AA7 AA8 AA9 AB10 AB11 AB12 AB13 AB14 AB15 AB16 AB17 AB18 AB19 AB2 AB20 AB21 AB22 AB23 AB4 AB5 AB6 AB7 AB8 AB9 AC1 AC10 AC11 AC13 AC14 AC16 AC17 AC19 AC2 AC20 AC22 AC23 AC4 AC5 AC7 AC8 B1 B10 B11 B12 B13 B14 B15 B16 B17 B18 B19 B2 B20 B21 B22 B23 B3 B4 B5 B6 B7 B8 B9 C10 C11 C12 C13 C14 C16 C17 C18 C19 C2 C20 C22 C3 C4 C5 C6 C7 C8 C9 D1 D10 D11 D13 D14 D16 D17 D19 D2 D20 D21 D22 D23 D3 D5 D7 D8 E1 E10 E11 E13 E14 E16 E17 E19 E2 E20 E21 E22 E23 E3 E4 E5 E7 E8 F12 F16 F17 F2 F21 F22 F3 F7 G1 G11 G13 G14 G16 G18 G19 G2 G20 G21 G22 G23 G3 G4 G5 G6 G7 G8 G9 H1 H13 H14 H15 H16 H19 H2 H20 H22 H23 H3 H4 H5 H6 J10 J11 J12 J13 J14 J15 J16 J2 J21 J3 J8 J9 K1 K10 K11 K12 K13 K14 K16 K18 K19 K2 K20 K22 K23 K3 K4 K5 K6 K7 K8 K9 L1 L10 L11 L12 L13 L14 L15 L16 L19 L2 L20 L22 L23 L3 L4 L5 L6 L7 L8 L9 M10 M11 M12 M13 M14 M15 M16 M2 M21 M22 M3 M4 M8 M9 N1 N10 N11 N12 N13 N14 N15 N16 N18 N19 N2 N20 N22 N23 N3 N4 N5 N6 N7 N8 N9 P1 P10 P11 P12 P13 P14 P16 P18 P19 P2 P20 P22 P23 P3 P5 P6 P7 P8 P9 R10 R11 R12 R13 R14 R15 R16 R2 R21 R22 R3 R4 R5 R6 R7 R8 R9 T1 T10 T11 T12 T13 T14 T15 T17 T19 T2 T20 T21 T22 T23 T3 T4 T6 T8 T9 U1 U11 U12 U15 U16 U18 U19 U2 U20 U21 U22 U23 U4 U5 U6 U7 U8 U9 V10 V14 V17 V18 V2 V21 V22 V3 V4 V5 V6 V8 V9 W1 W10 W11 W13 W16 W17 W19 W20 W21 W22 W23 W3 W4 W5 W7 W8 W9 Y10 Y11 Y13 Y14 Y16 Y17 Y19 Y2 Y21 Y22 Y23 Y3 Y4 Y6 Y7 Y8
* Stub for AllWinner-A64(FBGA396)
.ends

.subckt L 1 2
* Stub for L
.ends

.subckt MICRO_SD(TFC-WPAPR-08) 1 10 11 12 13 2 3 4 5 6 7 8 9
* Stub for MICRO_SD(TFC-WPAPR-08)
.ends

.subckt RA1206_(4x0603)_4B8_Smashed 1.1 1.2 2.1 2.2 3.1 3.2 4.1 4.2
* Stub for RA1206_(4x0603)_4B8_Smashed
.ends

.subckt AUDIO_JACK(SCJ325P00XG0B02G) 1 2 3 4 5
* Stub for AUDIO_JACK(SCJ325P00XG0B02G)
.ends

.subckt W25Q16BV 1 2 3 4 5 6 7 8
* Stub for W25Q16BV
.ends

.subckt SJ2W_Closed(1-2) 1 2 3
* Stub for SJ2W_Closed(1-2)
.ends

.subckt TESTPAD 1
* Stub for TESTPAD
.ends

.subckt Mounting_hole 0
* Stub for Mounting_hole
.ends

.subckt KLMAG2GEND-B031(FBGA153) A3 A4 A5 A6 B2 B3 B4 B5 B6 C2 C4 C6 E6 E7 F5 G5 H10 H5 J10 J5 K5 K8 K9 M4 M5 M6 N2 N4 N5 P3 P4 P5 P6
* Stub for KLMAG2GEND-B031(FBGA153)
.ends

.subckt SJ 1 2
* Stub for SJ
.ends

.subckt HDMI-SWM-19 0 1 10 11 12 13 14 15 16 17 18 19 2 3 4 5 6 7 8 9
* Stub for HDMI-SWM-19
.ends

.subckt RCLAMP0524P 1 10 2 3 4 5 6 7 8 9
* Stub for RCLAMP0524P
.ends

.subckt N-MOS+DIOD_Small 1 2 3
* Stub for N-MOS+DIOD_Small
.ends

.subckt USB-MINI 0 1 2 3 4 5
* Stub for USB-MINI
.ends

.subckt SY6280AAC(SOT23-5) 1 2 3 4 5
* Stub for SY6280AAC(SOT23-5)
.ends

.subckt RTL8723BS(ComboModule) 1 10 11 12 13 14 15 16 17 18 19 2 20 21 22 23 24 25 26 27 28 29 3 30 31 32 33 34 35 36 37 38 39 4 40 41 42 43 44 5 6 7 8 9
* Stub for RTL8723BS(ComboModule)
.ends

.subckt WIFI_ANT_ESP8266 1 2
* Stub for WIFI_ANT_ESP8266
.ends

.subckt LCD-ML40YA-V36P-2X20-LF 0 1 10 11 12 13 14 15 16 17 18 19 2 20 21 22 23 24 25 26 27 28 29 3 30 31 32 33 34 35 36 37 38 39 4 40 5 6 7 8 9
* Stub for LCD-ML40YA-V36P-2X20-LF
.ends

.subckt USB_A_VERTICAL 0 1 2 3 4
* Stub for USB_A_VERTICAL
.ends

.subckt KSZ9031RNXCC(QFN48_1DRILL(PADPITCH-0.5MM)) 1 10 11 12 13 14 15 16 17 18 19 2 20 21 22 23 24 25 26 27 28 29 3 30 31 32 33 34 35 36 37 38 39 4 40 41 42 43 44 45 46 47 48 49 5 6 7 8 9
* Stub for KSZ9031RNXCC(QFN48_1DRILL(PADPITCH-0.5MM))
.ends

.subckt TM211Q01FM22 1 10 11 12 13 14 2 3 4 5 6 7 8 9 SH1 SH2
* Stub for TM211Q01FM22
.ends

.subckt AMS1117-ADJ 1 2 3
* Stub for AMS1117-ADJ
.ends

.subckt JP1E 1 2
* Stub for JP1E
.ends

.subckt D 1 2
* Stub for D
.ends

.subckt AT24C16BN-SH(SO-8_150mil) 1 2 3 4 5 6 7 8
* Stub for AT24C16BN-SH(SO-8_150mil)
.ends

.subckt Crystal_GND 1 2 3
* Stub for Crystal_GND
.ends

.subckt D_Schottky 1 2
* Stub for D_Schottky
.ends

.subckt ESDS314DBVR(SOT-23-5) 1 2 3 4 5
* Stub for ESDS314DBVR(SOT-23-5)
.ends

.subckt AXP803 1 10 11 12 13 14 15 16 17 18 19 2 20 21 22 23 24 25 26 27 28 29 3 30 31 32 33 34 35 36 37 38 39 4 40 41 42 43 44 45 46 47 48 49 5 50 51 52 53 54 55 56 57 58 59 6 60 61 62 63 64 65 66 67 68 69 7 8 9
* Stub for AXP803
.ends

.subckt PWR-JAKPWR_JACK_UNI_MILLING + -
* Stub for PWR-JAKPWR_JACK_UNI_MILLING
.ends

.subckt FSMD035 1 2
* Stub for FSMD035
.ends

.subckt WPM1481 1 2 3 4 5 6 7 8
* Stub for WPM1481
.ends

.subckt LED 1 2
* Stub for LED
.ends

.subckt T1107A(6x3,8x2,5MM) 1 2
* Stub for T1107A(6x3,8x2,5MM)
.ends

.subckt Crystal 1 2
* Stub for Crystal
.ends

.subckt CON3 1 2 3
* Stub for CON3
.ends

.subckt BH10S 1 10 2 3 4 5 6 7 8 9
* Stub for BH10S
.ends

.subckt SMBJ6.0A 1 2
* Stub for SMBJ6.0A
.ends

.subckt CON2 1 2
* Stub for CON2
.ends

.subckt ML40YA-V36P-2X20-LF 1 10 11 12 13 14 15 16 17 18 19 2 20 21 22 23 24 25 26 27 28 29 3 30 31 32 33 34 35 36 37 38 39 4 40 5 6 7 8 9
* Stub for ML40YA-V36P-2X20-LF
.ends

.subckt GPH127SMT-02X10(PA-V16X-2X10-LF) 1 10 11 12 13 14 15 16 17 18 19 2 20 3 4 5 6 7 8 9
* Stub for GPH127SMT-02X10(PA-V16X-2X10-LF)
.ends

.subckt CON4 1 2 3 4
* Stub for CON4
.ends

.subckt SJ2W 1 2 3
* Stub for SJ2W
.ends

.subckt VDA2710NTA(SOT-23) 1 2 3
* Stub for VDA2710NTA(SOT-23)
.ends

.subckt P-MOS+DIOD 1 2 3
* Stub for P-MOS+DIOD
.ends

.subckt MT3608(SOT23-6) 1 2 3 4 5 6
* Stub for MT3608(SOT23-6)
.ends

