* Spice Netlist (renamed)

*--- Top Level ---
.subckt HDMI2USB DDR3_DDR0_A0 DDR3_DDR0_A1 DDR3_DDR0_A10 DDR3_DDR0_A11 DDR3_DDR0_A12 DDR3_DDR0_A13 DDR3_DDR0_A14 DDR3_DDR0_A2 DDR3_DDR0_A3 DDR3_DDR0_A4 DDR3_DDR0_A5 DDR3_DDR0_A6 DDR3_DDR0_A7 DDR3_DDR0_A8 DDR3_DDR0_A9 DDR3_DDR0_BA0 DDR3_DDR0_BA1 DDR3_DDR0_BA2 DDR3_DDR0_CAS_N DDR3_DDR0_CKE DDR3_DDR0_CK_N DDR3_DDR0_CK_P DDR3_DDR0_DQ0 DDR3_DDR0_DQ1 DDR3_DDR0_DQ10 DDR3_DDR0_DQ11 DDR3_DDR0_DQ12 DDR3_DDR0_DQ13 DDR3_DDR0_DQ14 DDR3_DDR0_DQ15 DDR3_DDR0_DQ2 DDR3_DDR0_DQ3 DDR3_DDR0_DQ4 DDR3_DDR0_DQ5 DDR3_DDR0_DQ6 DDR3_DDR0_DQ7 DDR3_DDR0_DQ8 DDR3_DDR0_DQ9 DDR3_DDR0_LDM DDR3_DDR0_LDQS_N DDR3_DDR0_LDQS_P DDR3_DDR0_ODT DDR3_DDR0_RAS_N DDR3_DDR0_RESET_N DDR3_DDR0_UDM DDR3_DDR0_UDQS_N DDR3_DDR0_UDQS_P DDR3_DDR0_WE_N DisplayPort_DPRXAUXCH_N DisplayPort_DPRXAUXCH_P DisplayPort_DPRXCONFIG1 DisplayPort_DPRXCONFIG2 DisplayPort_DPRX_LANEN0 DisplayPort_DPRX_LANEN1 DisplayPort_DPRX_LANEN2 DisplayPort_DPRX_LANEN3 DisplayPort_DPRX_LANEP0 DisplayPort_DPRX_LANEP1 DisplayPort_DPRX_LANEP2 DisplayPort_DPRX_LANEP3 DisplayPort_DPTXAUXCH_N DisplayPort_DPTXAUXCH_P DisplayPort_DPTXCONFIG1 DisplayPort_DPTXCONFIG2 DisplayPort_DPTX_LANEN0 DisplayPort_DPTX_LANEN1 DisplayPort_DPTX_LANEN2 DisplayPort_DPTX_LANEN3 DisplayPort_DPTX_LANEP0 DisplayPort_DPTX_LANEP1 DisplayPort_DPTX_LANEP2 DisplayPort_DPTX_LANEP3 Ethernet_AVDD3V3 Ethernet_ETH_INT_B Ethernet_ETH_MDC Ethernet_ETH_MDIO Ethernet_ETH_RESET_B Ethernet_ETH_RXCLK Ethernet_ETH_RXCTL Ethernet_ETH_RXD0 Ethernet_ETH_RXD1 Ethernet_ETH_RXD2 Ethernet_ETH_RXD3 Ethernet_ETH_TXCLK Ethernet_ETH_TXCTL Ethernet_ETH_TXD0 Ethernet_ETH_TXD1 Ethernet_ETH_TXD2 Ethernet_ETH_TXD3 Ethernet_ETH_VCC1V0 Ethernet_ETH_VCC3V3 Ethernet_LED0 Ethernet_LED1 Ethernet_MAC_SCL Ethernet_MAC_SDA Ethernet_MAC_WP Ethernet_VCC1V0 Ethernet_XTAL1_50MHZ Ethernet_XTAL2_50MHZ FPGA_Bank_0_3_DEBUG_IO0 FPGA_Bank_0_3_DEBUG_IO1 FPGA_Bank_0_3_DIFFCLK_A0N FPGA_Bank_0_3_DIFFCLK_A0P FPGA_Bank_0_3_DIFFCLK_A1N FPGA_Bank_0_3_DIFFCLK_A1P FPGA_Bank_0_3_DIFFCLK_B0N FPGA_Bank_0_3_DIFFCLK_B0P FPGA_Bank_0_3_DIFFCLK_B1N FPGA_Bank_0_3_DIFFCLK_B1P FPGA_Bank_0_3_DIFFCLK_XN FPGA_Bank_0_3_DIFFCLK_XP FPGA_Bank_0_3_DIFFIO_A0N FPGA_Bank_0_3_DIFFIO_A0P FPGA_Bank_0_3_DIFFIO_A1N FPGA_Bank_0_3_DIFFIO_A1P FPGA_Bank_0_3_DIFFIO_A2N FPGA_Bank_0_3_DIFFIO_A2P FPGA_Bank_0_3_DIFFIO_A3N FPGA_Bank_0_3_DIFFIO_A3P FPGA_Bank_0_3_DIFFIO_A4N FPGA_Bank_0_3_DIFFIO_A4P FPGA_Bank_0_3_DIFFIO_A5N FPGA_Bank_0_3_DIFFIO_A5P FPGA_Bank_0_3_DIFFIO_A6N FPGA_Bank_0_3_DIFFIO_A6P FPGA_Bank_0_3_DIFFIO_B0N FPGA_Bank_0_3_DIFFIO_B0P FPGA_Bank_0_3_DIFFIO_B1N FPGA_Bank_0_3_DIFFIO_B1P FPGA_Bank_0_3_DIFFIO_B2N FPGA_Bank_0_3_DIFFIO_B2P FPGA_Bank_0_3_DIFFIO_B3N FPGA_Bank_0_3_DIFFIO_B3P FPGA_Bank_0_3_DIFFIO_B4N FPGA_Bank_0_3_DIFFIO_B4P FPGA_Bank_0_3_DIFFIO_B5N FPGA_Bank_0_3_DIFFIO_B5P FPGA_Bank_0_3_DIFFIO_B6N FPGA_Bank_0_3_DIFFIO_B6P FPGA_Bank_0_3_DIFFIO_XN FPGA_Bank_0_3_DIFFIO_XP FPGA_Bank_0_3_DIFFIO_YN FPGA_Bank_0_3_DIFFIO_YP FPGA_Bank_0_3_DIFFIO_ZN FPGA_Bank_0_3_DIFFIO_ZP FPGA_Bank_0_3_HSWAP FPGA_Bank_0_3_MGT135MHz_N FPGA_Bank_0_3_MGT135MHz_P FPGA_Bank_0_3_MGTREFCLK0_101_N FPGA_Bank_0_3_MGTREFCLK0_101_P FPGA_Bank_0_3_MGTSMACLK_N FPGA_Bank_0_3_MGTSMACLK_P FPGA_Bank_0_3_PCIE_RESET FPGA_Bank_0_3_PCIO0 FPGA_Bank_0_3_PCIO1 FPGA_Bank_0_3_PCIO2 FPGA_Bank_0_3_PCIO3 FPGA_Bank_0_3_SMCLK FPGA_Bank_0_3_SMDATA FPGA_Bank_0_3_SWITCH FPGA_Bank_1_2_100MHz FPGA_Bank_1_2_CYPRESS_RESET FPGA_Bank_1_2_CY_CTL0 FPGA_Bank_1_2_CY_CTL1 FPGA_Bank_1_2_CY_CTL2 FPGA_Bank_1_2_CY_CTL3 FPGA_Bank_1_2_CY_CTL4 FPGA_Bank_1_2_CY_CTL5 FPGA_Bank_1_2_CY_FD0 FPGA_Bank_1_2_CY_FD1 FPGA_Bank_1_2_CY_FD10 FPGA_Bank_1_2_CY_FD11 FPGA_Bank_1_2_CY_FD12 FPGA_Bank_1_2_CY_FD13 FPGA_Bank_1_2_CY_FD14 FPGA_Bank_1_2_CY_FD15 FPGA_Bank_1_2_CY_FD2 FPGA_Bank_1_2_CY_FD3 FPGA_Bank_1_2_CY_FD4 FPGA_Bank_1_2_CY_FD5 FPGA_Bank_1_2_CY_FD6 FPGA_Bank_1_2_CY_FD7 FPGA_Bank_1_2_CY_FD8 FPGA_Bank_1_2_CY_FD9 FPGA_Bank_1_2_CY_IFCLK FPGA_Bank_1_2_CY_INT5 FPGA_Bank_1_2_CY_PA0 FPGA_Bank_1_2_CY_PA1 FPGA_Bank_1_2_CY_PA2 FPGA_Bank_1_2_CY_PA3 FPGA_Bank_1_2_CY_PA4 FPGA_Bank_1_2_CY_PA5 FPGA_Bank_1_2_CY_PA6 FPGA_Bank_1_2_CY_PA7 FPGA_Bank_1_2_CY_PC0 FPGA_Bank_1_2_CY_PC1 FPGA_Bank_1_2_CY_PC2 FPGA_Bank_1_2_CY_PC3 FPGA_Bank_1_2_CY_PC4 FPGA_Bank_1_2_CY_PC5 FPGA_Bank_1_2_CY_PC6 FPGA_Bank_1_2_CY_PC7 FPGA_Bank_1_2_CY_RD FPGA_Bank_1_2_CY_RD0 FPGA_Bank_1_2_CY_RD1 FPGA_Bank_1_2_CY_RD2 FPGA_Bank_1_2_CY_RD3 FPGA_Bank_1_2_CY_RD4 FPGA_Bank_1_2_CY_RD5 FPGA_Bank_1_2_CY_RXD0 FPGA_Bank_1_2_CY_RXD1 FPGA_Bank_1_2_CY_T0 FPGA_Bank_1_2_CY_TXD0 FPGA_Bank_1_2_CY_TXD1 FPGA_Bank_1_2_CY_WR FPGA_Bank_1_2_DPRXHPD FPGA_Bank_1_2_DPTXHPD FPGA_Bank_1_2_FPGA_M0_CMP_MISO FPGA_Bank_1_2_FPGA_M1 FPGA_Bank_1_2_INIT_B FPGA_Bank_1_2_SD_CLK FPGA_Bank_1_2_SD_CMD FPGA_Bank_1_2_SD_DAT0 FPGA_Bank_1_2_SD_DAT1 FPGA_Bank_1_2_SD_DAT2 FPGA_Bank_1_2_SD_DAT3 FPGA_Bank_1_2_SPI_CLK FPGA_Bank_1_2_SPI_CS_N FPGA_Bank_1_2_SPI_D1_MISO2 FPGA_Bank_1_2_SPI_D2_MISO3 FPGA_Bank_1_2_SPI_DO_DIN_MISO1 FPGA_Bank_1_2_SPI_MOSI_CSI_N_MISO0 FPGA_Bank_1_2_TMDS_RX1_0_N FPGA_Bank_1_2_TMDS_RX1_0_P FPGA_Bank_1_2_TMDS_RX1_1_N FPGA_Bank_1_2_TMDS_RX1_1_P FPGA_Bank_1_2_TMDS_RX1_2_N FPGA_Bank_1_2_TMDS_RX1_2_P FPGA_Bank_1_2_TMDS_RX1_CEC FPGA_Bank_1_2_TMDS_RX1_CLK_N FPGA_Bank_1_2_TMDS_RX1_CLK_P FPGA_Bank_1_2_TMDS_RX1_HOT FPGA_Bank_1_2_TMDS_RX1_SCL FPGA_Bank_1_2_TMDS_RX1_SDA FPGA_Bank_1_2_TMDS_RX2_0_N FPGA_Bank_1_2_TMDS_RX2_0_P FPGA_Bank_1_2_TMDS_RX2_1_N FPGA_Bank_1_2_TMDS_RX2_1_P FPGA_Bank_1_2_TMDS_RX2_2_N FPGA_Bank_1_2_TMDS_RX2_2_P FPGA_Bank_1_2_TMDS_RX2_CEC FPGA_Bank_1_2_TMDS_RX2_CLK_N FPGA_Bank_1_2_TMDS_RX2_CLK_P FPGA_Bank_1_2_TMDS_RX2_HOT FPGA_Bank_1_2_TMDS_RX2_SCL FPGA_Bank_1_2_TMDS_RX2_SDA FPGA_Bank_1_2_TMDS_TX1_0_N FPGA_Bank_1_2_TMDS_TX1_0_P FPGA_Bank_1_2_TMDS_TX1_1_N FPGA_Bank_1_2_TMDS_TX1_1_P FPGA_Bank_1_2_TMDS_TX1_2_N FPGA_Bank_1_2_TMDS_TX1_2_P FPGA_Bank_1_2_TMDS_TX1_CEC FPGA_Bank_1_2_TMDS_TX1_CLK_N FPGA_Bank_1_2_TMDS_TX1_CLK_P FPGA_Bank_1_2_TMDS_TX1_HOT FPGA_Bank_1_2_TMDS_TX1_SCL FPGA_Bank_1_2_TMDS_TX1_SDA FPGA_Bank_1_2_TMDS_TX2_0_N FPGA_Bank_1_2_TMDS_TX2_0_P FPGA_Bank_1_2_TMDS_TX2_1_N FPGA_Bank_1_2_TMDS_TX2_1_P FPGA_Bank_1_2_TMDS_TX2_2_N FPGA_Bank_1_2_TMDS_TX2_2_P FPGA_Bank_1_2_TMDS_TX2_CEC FPGA_Bank_1_2_TMDS_TX2_CLK_N FPGA_Bank_1_2_TMDS_TX2_CLK_P FPGA_Bank_1_2_TMDS_TX2_HOT FPGA_Bank_1_2_TMDS_TX2_SCL FPGA_Bank_1_2_TMDS_TX2_SDA FPGA_Bank_1_2_USB_D0 FPGA_Bank_1_2_USB_D1 FPGA_Bank_1_2_USB_D2 FPGA_Bank_1_2_USB_D3 FPGA_Bank_1_2_USB_D4 FPGA_Bank_1_2_USB_D5 FPGA_Bank_1_2_USB_D6 FPGA_Bank_1_2_USB_D7 FPGA_Bank_1_2_USB_DIR FPGA_Bank_1_2_USB_NXT FPGA_Bank_1_2_USB_REFCLK FPGA_Bank_1_2_USB_RESETB FPGA_Bank_1_2_USB_STP FPGA_Power_DONE FPGA_Power_PROG_B FPGA_Power_RFS FPGA_Power_SUSPEND FPGA_Power_TCK FPGA_Power_TMS FPGA_Power_VBATT FPGA_Power_VFS GND GPIOs_PRSNT HDMI_HDMI_TX1_VCC5V0 HDMI_HDMI_TX2_VCC5V0 HDMI_HDMI_VCC5V0 HDMI_P1_CEC HDMI_P1_HOT HDMI_P1_SCL HDMI_P1_SDA HDMI_P2_CEC HDMI_P2_HOT HDMI_P2_SCL HDMI_P2_SDA HDMI_P3_CEC HDMI_P3_HOT HDMI_P3_SCL HDMI_P3_SDA HDMI_P4_CEC HDMI_P4_HOT HDMI_P4_SCL HDMI_P4_SDA Power_Conference_12V Power_Consumer_12V Power_VIN_48 Power_VIN__48V Power_VIN__48V_0 SPI_Flash_27MHz SPI_Flash_RST SPI_Flash_TDO_FPGA_TDO_JTAG SPI_Flash_TDO_USB_TDI_FPGA USB_CPEN USB_CYDN USB_CYDP USB_CYP_RESET USB_ID USB_U1_SDA USB_USB_5V USB_USB_DM USB_USB_DP USB_XTALIN USB_XTALIOUT VCC12V0 VCC1V2 VCC1V5 VCC3V3 VCC4V0 VTTDDR0 VTTREF unnamed
  XU8 VCC1V5 unnamed unnamed unnamed VCC12V0 VCC12V0 GND unnamed unnamed unnamed GND unnamed unnamed GND GND TPS54625
  XC150 unnamed unnamed C
  XL4 unnamed VCC1V5 INDUCTOR
  XR112 VCC1V5 unnamed R
  XR113 unnamed GND R
  XC143 GND unnamed C
  XR102 unnamed unnamed R
  XC137 GND unnamed C
  XR100 VCC12V0 unnamed R
  XC133 GND VCC12V0 C
  XC79 GND VCC12V0 C
  XC161 GND VCC1V5 C
  XU9 VCC1V2 unnamed unnamed unnamed VCC12V0 VCC12V0 GND unnamed unnamed unnamed GND unnamed unnamed GND GND TPS54625
  XC152 unnamed unnamed C
  XL5 unnamed VCC1V2 INDUCTOR
  XR114 VCC1V2 unnamed R
  XR115 unnamed GND R
  XC144 GND unnamed C
  XR104 unnamed unnamed R
  XC141 GND unnamed C
  XR103 VCC12V0 unnamed R
  XC140 GND VCC12V0 C
  XC134 GND VCC12V0 C
  XC164 GND VCC1V2 C
  XU7 unnamed unnamed unnamed VCC12V0 VCC12V0 VCC12V0 VCC12V0 VCC12V0 VCC12V0 unnamed VCC12V0 unnamed unnamed unnamed unnamed GND unnamed unnamed unnamed unnamed unnamed unnamed unnamed TPS53319
  XR107 GND unnamed R
  XC148 GND unnamed C
  XR108 unnamed unnamed R
  XC149 unnamed unnamed C
  XR98 unnamed GND R
  XR95 VCC12V0 unnamed R
  XR96 unnamed GND R
  XR97 unnamed unnamed R
  XC77 GND VCC12V0 C
  XC75 GND VCC12V0 C
  XC72 GND VCC12V0 C
  XL3 unnamed VCC4V0 INDUCTOR
  XR109 unnamed unnamed R
  XC154 VCC4V0 unnamed C
  XC151 unnamed unnamed C
  XR110 unnamed VCC4V0 R
  XR111 GND unnamed R
  XC157 GND VCC4V0 C
  XC59 GND Power_Consumer_12V C
  XC61 GND Power_Consumer_12V C
  XR101 VCC1V5 unnamed R
  XR105 unnamed GND R
  XC146 unnamed GND C
  XC81 GND VCC1V5 C
  XC138 GND VCC1V5 C
  XC156 GND VTTDDR0 C
  XC159 GND VTTDDR0 C
  XC162 GND VTTDDR0 C
  XR106 unnamed VCC3V3 R
  XC147 GND VCC3V3 C
  XC153 GND VTTREF C
  XC73 GND VCC12V0 C
  XC74 GND VCC12V0 C
  XC78 VCC12V0 GND C
  XC135 VCC12V0 GND C
  XC165 GND VCC1V5 C
  XC160 GND VCC4V0 C
  XC163 GND VCC4V0 C
  XC136 VCC1V5 GND C
  XC76 GND VCC1V5 C
  XC166 GND VTTDDR0 C
  XC168 GND VTTDDR0 C
  XC167 GND VCC1V2 C
  XC139 GND VCC12V0 C
  XC145 GND VCC12V0 C
  XR99 unnamed GND R
  XC155 unnamed VCC1V5 C
  XC142 VCC12V0 GND C
  XC158 VCC1V2 unnamed C
  XC80 VCC12V0 GND C
  XP1 Power_VIN__48V Power_VIN__48V_0 CONN_2
  XU6 unnamed Power_VIN_48 unnamed unnamed unnamed unnamed GND unnamed GND TPS54560
  XU4 Power_VIN_48 Power_VIN__48V_0 Power_VIN__48V GND GBU15005-G
  XC60 unnamed unnamed C
  XR90 unnamed Power_Conference_12V R
  XD5 GND unnamed DIODE
  XC57 GND Power_VIN_48 C
  XC56 GND Power_VIN_48 C
  XC55 GND Power_VIN_48 C
  XR77 unnamed Power_VIN_48 R
  XR78 unnamed GND R
  XR79 unnamed GND R
  XL2 unnamed Power_Conference_12V INDUCTOR
  XR91 GND unnamed R
  XC67 GND Power_Conference_12V C
  XC68 GND Power_Conference_12V C
  XC69 GND Power_Conference_12V C
  XC51 GND Power_VIN_48 C
  XC63 unnamed GND C
  XR87 unnamed unnamed R
  XC65 GND unnamed C
  XC70 GND Power_Conference_12V C
  XC71 GND Power_Conference_12V C
  XC48 GND Power_VIN_48 C
  XC45 GND Power_VIN_48 C
  XCON1 Power_VIN__48V_0 Power_VIN__48V Power_VIN__48V BARREL_JACK
  XCON2 Power_Consumer_12V GND GND BARREL_JACK
  XD6 Power_Conference_12V unnamed DIODESCH
  XD9 Power_Consumer_12V unnamed DIODESCH
  XD8 Power_Consumer_12V unnamed DIODESCH
  XD7 Power_Conference_12V unnamed DIODESCH
  XF1 unnamed VCC12V0 FUSE
  XU12 unnamed VCC3V3 GND VCC1V5 VTTDDR0 GND VTTDDR0 VTTREF VCC3V3 GND unnamed TPS51200
  XD10 unnamed GND LED
  XR94 VCC12V0 unnamed R
  XD4 VCC4V0 VCC3V3 DIODE
  XP27 unnamed unnamed unnamed GND GND GND ATX_POWER_SUPPLY
  XD14 unnamed VCC12V0 DIODESCH
  XC268 GND VCC12V0 C
  XC269 GND VCC12V0 C
  XU10 GND unnamed GND unnamed GND DisplayPort_DPTX_LANEN2 VCC1V2 DisplayPort_DPTX_LANEN3 FPGA_Bank_0_3_DIFFIO_B2N FPGA_Bank_0_3_DIFFIO_A1N FPGA_Bank_0_3_DIFFIO_XN FPGA_Bank_0_3_DIFFIO_A6N FPGA_Bank_0_3_DIFFIO_B0N FPGA_Power_TCK GND FPGA_Bank_0_3_DIFFIO_B6N FPGA_Bank_0_3_DIFFIO_A5N FPGA_Bank_0_3_DIFFIO_B5N DisplayPort_DPTX_LANEN0 VCC1V2 DisplayPort_DPTX_LANEN1 GND FPGA_Bank_0_3_DEBUG_IO1 FPGA_Bank_1_2_TMDS_TX1_1_P VCC3V3 Ethernet_ETH_RXCLK GND FPGA_Bank_1_2_USB_D4 VCC3V3 FPGA_Bank_1_2_TMDS_TX2_1_P GND FPGA_Bank_1_2_TMDS_TX2_CEC VCC3V3 FPGA_Bank_0_3_DEBUG_IO0 FPGA_Bank_1_2_SPI_DO_DIN_MISO1 FPGA_Bank_1_2_FPGA_M0_CMP_MISO FPGA_Power_SUSPEND FPGA_Bank_1_2_SPI_CS_N FPGA_Bank_1_2_SD_DAT0 GND Ethernet_ETH_TXD2 VCC3V3 DisplayPort_DPRXCONFIG1 GND GND FPGA_Bank_1_2_TMDS_TX1_1_N FPGA_Bank_1_2_TMDS_TX1_CLK_N Ethernet_ETH_TXCLK FPGA_Bank_1_2_100MHz FPGA_Bank_1_2_USB_D5 FPGA_Bank_1_2_TMDS_TX2_0_N FPGA_Bank_1_2_TMDS_TX2_1_N FPGA_Bank_1_2_TMDS_TX2_SDA FPGA_Bank_1_2_TMDS_TX2_HOT DisplayPort_DPTXCONFIG2 FPGA_Power_PROG_B FPGA_Bank_1_2_SPI_MOSI_CSI_N_MISO0 FPGA_Power_DONE GND VCC3V3 FPGA_Bank_1_2_SD_DAT1 FPGA_Bank_1_2_SD_DAT2 Ethernet_ETH_TXD3 FPGA_Bank_1_2_TMDS_TX1_HOT DisplayPort_DPRXCONFIG2 FPGA_Bank_1_2_TMDS_TX1_2_N VTTREF unnamed GND unnamed VCC1V2 DisplayPort_DPTX_LANEP2 GND DisplayPort_DPTX_LANEP3 GND FPGA_Bank_0_3_DIFFIO_A1P VCC3V3 FPGA_Bank_0_3_DIFFIO_A6P FPGA_Bank_0_3_DIFFIO_B0P FPGA_Bank_1_2_CY_PA4 FPGA_Bank_1_2_CY_PA5 FPGA_Bank_0_3_DIFFIO_B6P VCC3V3 GND DisplayPort_DPTX_LANEP0 GND DisplayPort_DPTX_LANEP1 VCC1V2 Ethernet_MAC_SDA VCC1V2 FPGA_Bank_0_3_MGTSMACLK_P GND DisplayPort_DPRX_LANEN1 GND DisplayPort_DPRX_LANEN0 GND FPGA_Bank_0_3_DIFFIO_B2P FPGA_Bank_0_3_DIFFIO_A0N FPGA_Bank_0_3_DIFFIO_XP VCC1V5 FPGA_Bank_1_2_CY_FD0 VCC3V3 FPGA_Bank_1_2_CY_FD1 FPGA_Bank_0_3_HSWAP FPGA_Bank_0_3_DIFFIO_A5P FPGA_Bank_0_3_DIFFIO_B5P GND DisplayPort_DPRX_LANEN3 GND DisplayPort_DPRX_LANEN2 unnamed GND FPGA_Bank_0_3_MGTSMACLK_N VCC1V2 DisplayPort_DPRX_LANEP1 VCC1V2 DisplayPort_DPRX_LANEP0 GND FPGA_Bank_0_3_DIFFIO_A0P FPGA_Bank_0_3_DIFFCLK_XP FPGA_Bank_0_3_DIFFCLK_XN unnamed FPGA_Power_TMS FPGA_Bank_1_2_CY_FD4 FPGA_Bank_1_2_CY_FD5 FPGA_Bank_0_3_PCIE_RESET FPGA_Bank_0_3_DIFFIO_B4P FPGA_Bank_0_3_DIFFIO_B4N GND DisplayPort_DPRX_LANEP3 VCC1V2 DisplayPort_DPRX_LANEP2 DDR3_DDR0_A11 VCC1V2 GND FPGA_Bank_0_3_MGT135MHz_P VCC1V2 GND GND FPGA_Bank_0_3_DIFFCLK_B0N VCC3V3 SPI_Flash_TDO_USB_TDI_FPGA VCC3V3 GND FPGA_Bank_1_2_CY_FD12 GND FPGA_Bank_1_2_CY_FD13 DDR3_DDR0_RESET_N unnamed FPGA_Bank_0_3_DIFFIO_A4P FPGA_Bank_0_3_DIFFIO_A4N GND VCC1V2 unnamed DDR3_DDR0_A12 FPGA_Bank_0_3_DIFFCLK_A1P VCC3V3 FPGA_Bank_0_3_MGT135MHz_N GND FPGA_Bank_0_3_DIFFCLK_A0P FPGA_Bank_0_3_DIFFCLK_A0N FPGA_Bank_0_3_DIFFCLK_B0P FPGA_Bank_0_3_DIFFIO_B1N FPGA_Bank_1_2_CY_PA0 FPGA_Bank_1_2_CY_PA1 DDR3_DDR0_CKE FPGA_Bank_1_2_CY_FD7 FPGA_Bank_1_2_CY_FD10 FPGA_Bank_1_2_CY_FD11 unnamed VCC1V5 FPGA_Bank_0_3_PCIO3 VCC3V3 FPGA_Bank_0_3_DIFFIO_YP FPGA_Bank_0_3_DIFFIO_YN FPGA_Bank_0_3_DIFFIO_ZN DDR3_DDR0_A9 VCC3V3 FPGA_Bank_0_3_DIFFCLK_B1N VCC3V3 FPGA_Bank_0_3_DIFFIO_A3N VCC3V3 FPGA_Bank_0_3_DIFFIO_A2N FPGA_Bank_0_3_DIFFIO_B1P SPI_Flash_TDO_FPGA_TDO_JTAG GND FPGA_Bank_1_2_CY_FD6 VCC1V5 FPGA_Bank_1_2_CY_T0 VCC3V3 FPGA_Bank_1_2_CYPRESS_RESET DDR3_DDR0_A8 unnamed GND Ethernet_MAC_SCL FPGA_Bank_0_3_PCIO0 FPGA_Bank_0_3_DIFFIO_ZP FPGA_Bank_0_3_DIFFCLK_A1N DDR3_DDR0_BA2 FPGA_Bank_0_3_DIFFIO_B3P FPGA_Bank_0_3_DIFFIO_B3N FPGA_Bank_0_3_DIFFCLK_B1P FPGA_Bank_0_3_DIFFIO_A3P FPGA_Bank_0_3_DIFFIO_A2P VCC3V3 FPGA_Bank_1_2_CY_PA2 FPGA_Bank_1_2_CY_PA3 FPGA_Bank_1_2_CY_FD8 FPGA_Bank_1_2_CY_FD9 DDR3_DDR0_WE_N FPGA_Bank_1_2_CY_FD15 FPGA_Bank_1_2_TMDS_RX1_1_P FPGA_Bank_1_2_TMDS_RX1_1_N DDR3_DDR0_A4 unnamed DDR3_DDR0_A14 unnamed GND FPGA_Bank_0_3_PCIO2 VCC3V3 DDR3_DDR0_BA1 VCC1V2 GND VCC1V2 GND VCC1V2 GND FPGA_Bank_1_2_CY_PA6 FPGA_Bank_1_2_CY_PA7 VCC3V3 FPGA_Bank_1_2_CY_FD14 GND FPGA_Bank_1_2_TMDS_RX1_0_P GND FPGA_Bank_1_2_TMDS_RX1_0_N DDR3_DDR0_BA0 DDR3_DDR0_A10 VCC1V5 DDR3_DDR0_A13 FPGA_Bank_0_3_PCIO1 VCC1V2 GND DDR3_DDR0_A1 GND VCC1V2 GND VCC1V2 GND VCC3V3 FPGA_Bank_1_2_CY_FD3 FPGA_Bank_1_2_TMDS_RX1_CEC FPGA_Bank_1_2_CY_WR FPGA_Bank_1_2_CY_RD DDR3_DDR0_A0 FPGA_Bank_1_2_TMDS_RX1_2_P FPGA_Bank_0_3_MGTREFCLK0_101_P FPGA_Bank_0_3_MGTREFCLK0_101_N DDR3_DDR0_CK_N DDR3_DDR0_CK_P DDR3_DDR0_A2 DDR3_DDR0_A7 unnamed VTTREF VCC1V2 DDR3_DDR0_DQ5 VCC1V2 GND VCC1V2 GND VCC1V2 FPGA_Bank_1_2_CY_FD2 VCC3V3 FPGA_Bank_1_2_TMDS_RX1_SCL GND FPGA_Bank_1_2_TMDS_RX1_2_N VCC1V5 FPGA_Bank_1_2_TMDS_RX2_CLK_P VCC3V3 FPGA_Bank_1_2_TMDS_RX2_CLK_N DDR3_DDR0_DQ4 DDR3_DDR0_A6 GND DDR3_DDR0_ODT VCC1V5 VCC3V3 GND DDR3_DDR0_DQ7 GND VCC1V2 GND VCC1V2 GND VCC3V3 FPGA_Bank_1_2_CY_RD2 FPGA_Bank_1_2_CY_CTL4 FPGA_Bank_1_2_CY_CTL3 FPGA_Bank_1_2_TMDS_RX1_CLK_N DDR3_DDR0_DQ6 FPGA_Bank_1_2_TMDS_RX1_CLK_P FPGA_Bank_1_2_TMDS_RX2_0_P FPGA_Bank_1_2_TMDS_RX2_0_N DDR3_DDR0_A5 DDR3_DDR0_CAS_N DDR3_DDR0_RAS_N DDR3_DDR0_A3 unnamed VTTREF VCC1V2 DDR3_DDR0_LDQS_N VCC1V2 GND VCC1V2 GND VCC1V2 FPGA_Bank_1_2_CY_RD3 FPGA_Bank_1_2_CY_CTL0 GND VCC3V3 SPI_Flash_27MHz GND FPGA_Bank_1_2_TMDS_RX2_1_P GND FPGA_Bank_1_2_TMDS_RX2_1_N DDR3_DDR0_LDQS_P DDR3_DDR0_LDM VCC1V5 FPGA_Bank_0_3_SMCLK FPGA_Bank_0_3_SMDATA VCC3V3 GND DDR3_DDR0_DQ3 GND VCC1V2 GND VCC1V2 GND FPGA_Power_RFS FPGA_Bank_1_2_CY_CTL1 FPGA_Bank_1_2_CY_RXD1 FPGA_Bank_1_2_CY_RXD0 FPGA_Bank_1_2_CY_RD0 DDR3_DDR0_DQ2 FPGA_Bank_1_2_CY_IFCLK FPGA_Bank_1_2_TMDS_RX2_2_P FPGA_Bank_1_2_TMDS_RX2_2_N DDR3_DDR0_UDM unnamed unnamed unnamed unnamed VTTREF VCC1V2 DDR3_DDR0_DQ1 VCC3V3 DisplayPort_DPRXAUXCH_P VCC3V3 FPGA_Bank_1_2_SPI_D1_MISO2 VCC1V2 FPGA_Bank_1_2_CY_CTL2 FPGA_Bank_1_2_CY_CTL5 FPGA_Bank_1_2_CY_TXD1 GND FPGA_Bank_1_2_CY_RD1 VCC1V5 FPGA_Bank_1_2_TMDS_RX2_HOT VCC3V3 FPGA_Bank_1_2_TMDS_RX2_SDA DDR3_DDR0_DQ0 unnamed GND VCC3V3 unnamed Ethernet_ETH_RXD1 Ethernet_ETH_RXD0 DDR3_DDR0_DQ9 DisplayPort_DPRXAUXCH_P DisplayPort_DPRXAUXCH_N FPGA_Bank_1_2_TMDS_TX2_CLK_P VCC3V3 FPGA_Bank_1_2_SPI_D2_MISO3 DisplayPort_DPTXAUXCH_P FPGA_Power_VBATT FPGA_Bank_1_2_CY_TXD0 FPGA_Bank_1_2_TMDS_RX1_SDA FPGA_Bank_1_2_CY_INT5 DDR3_DDR0_DQ8 FPGA_Bank_1_2_CY_RD5 FPGA_Bank_1_2_TMDS_RX2_SCL FPGA_Bank_1_2_TMDS_RX2_CEC unnamed unnamed unnamed unnamed FPGA_Bank_1_2_SD_CLK Ethernet_ETH_MDIO VCC3V3 DDR3_DDR0_DQ11 DisplayPort_DPRXAUXCH_N VCC3V3 FPGA_Bank_1_2_TMDS_TX2_CLK_N FPGA_Bank_1_2_TMDS_TX2_2_N FPGA_Bank_1_2_TMDS_TX2_2_P DisplayPort_DPTXAUXCH_N DisplayPort_DPTXAUXCH_P FPGA_Power_VFS VCC3V3 FPGA_Bank_1_2_CY_RD4 GND FPGA_Bank_1_2_CY_PC0 GND FPGA_Bank_1_2_CY_PC1 DDR3_DDR0_DQ10 unnamed VCC1V5 FPGA_Bank_1_2_SD_CMD GND Ethernet_ETH_RESET_B Ethernet_ETH_RXCTL DDR3_DDR0_UDQS_N GND FPGA_Bank_1_2_DPTXHPD VCC3V3 FPGA_Bank_1_2_USB_NXT GND DisplayPort_DPTXAUXCH_N VCC3V3 FPGA_Bank_1_2_USB_RESETB unnamed FPGA_Bank_1_2_TMDS_RX1_HOT DDR3_DDR0_UDQS_P DisplayPort_DPTXCONFIG1 FPGA_Bank_1_2_CY_PC2 FPGA_Bank_1_2_CY_PC3 unnamed GND unnamed VCC3V3 Ethernet_ETH_MDC VCC3V3 Ethernet_ETH_INT_B DDR3_DDR0_DQ13 FPGA_Bank_1_2_TMDS_TX1_CEC FPGA_Bank_1_2_DPRXHPD FPGA_Bank_1_2_TMDS_TX1_0_P FPGA_Bank_1_2_USB_DIR FPGA_Bank_1_2_USB_D1 FPGA_Bank_1_2_USB_D7 GND FPGA_Bank_1_2_USB_D3 FPGA_Bank_1_2_USB_STP GND VCC1V5 FPGA_Bank_1_2_CY_PC4 VCC3V3 FPGA_Bank_1_2_CY_PC5 DDR3_DDR0_DQ12 unnamed VCC3V3 Ethernet_ETH_RXD2 GND Ethernet_ETH_TXCTL Ethernet_ETH_TXD0 DDR3_DDR0_DQ15 FPGA_Bank_1_2_TMDS_TX1_SDA FPGA_Bank_1_2_TMDS_TX1_CLK_P FPGA_Bank_1_2_TMDS_TX1_0_N FPGA_Bank_1_2_USB_REFCLK FPGA_Bank_1_2_USB_D0 FPGA_Bank_1_2_TMDS_TX2_0_P FPGA_Bank_1_2_USB_D6 FPGA_Bank_1_2_TMDS_TX2_SCL FPGA_Bank_1_2_USB_D2 FPGA_Bank_1_2_FPGA_M1 DDR3_DDR0_DQ14 FPGA_Bank_1_2_SPI_CLK FPGA_Bank_1_2_CY_PC6 FPGA_Bank_1_2_CY_PC7 FPGA_Bank_0_3_SWITCH FPGA_Bank_1_2_INIT_B FPGA_Bank_1_2_SD_DAT3 Ethernet_ETH_RXD3 FPGA_Bank_1_2_TMDS_TX1_SCL Ethernet_ETH_TXD1 FPGA_Bank_1_2_TMDS_TX1_2_P XC6SLX150T
  XR53 FPGA_Bank_0_3_HSWAP GND R
  XR57 FPGA_Power_RFS VCC3V3 R
  XC82 VCC1V5 GND C
  XC84 VCC1V5 GND C
  XC86 VCC1V5 GND C
  XC88 VCC1V5 GND C
  XC90 VCC1V2 GND C
  XC92 VCC1V5 GND C
  XC94 VCC1V5 GND C
  XC96 VCC1V5 GND C
  XC98 VCC1V5 GND C
  XC102 VCC1V5 GND C
  XC108 GND VCC3V3 C
  XC110 GND VCC3V3 C
  XC112 GND VCC3V3 C
  XC114 GND VCC3V3 C
  XC83 GND VCC3V3 C
  XC85 GND VCC3V3 C
  XC87 GND VCC3V3 C
  XC89 GND VCC3V3 C
  XC91 GND VCC3V3 C
  XC93 GND VCC3V3 C
  XC95 GND VCC3V3 C
  XC97 GND VCC3V3 C
  XC99 GND VCC3V3 C
  XC101 GND VCC3V3 C
  XC103 GND VCC3V3 C
  XC105 GND VCC3V3 C
  XC107 GND VCC3V3 C
  XC109 GND VCC3V3 C
  XC111 GND VCC3V3 C
  XC115 GND VCC3V3 C
  XC117 GND VCC3V3 C
  XC119 GND VCC3V3 C
  XC121 VCC1V2 GND C
  XC123 GND VCC3V3 C
  XC125 GND VCC3V3 C
  XC127 VCC1V5 GND C
  XC116 GND VCC3V3 C
  XC118 GND VCC3V3 C
  XC120 GND VCC3V3 C
  XC122 VCC1V2 GND C
  XC124 VCC1V2 GND C
  XC126 VCC1V2 GND C
  XC128 VCC1V2 GND C
  XC129 VCC1V2 GND C
  XC130 VCC1V2 GND C
  XC131 VCC1V2 GND C
  XD1 unnamed FPGA_Power_DONE LED
  XR55 unnamed VCC3V3 R
  XR56 FPGA_Power_PROG_B VCC3V3 R
  XR52 VCC3V3 FPGA_Bank_1_2_INIT_B R
  XC190 GND VCC3V3 C
  XC213 GND VCC3V3 C
  XC215 VCC1V2 GND C
  XC221 VCC1V2 GND C
  XC236 VCC1V2 GND C
  XC237 VCC1V2 GND C
  XR29 GND FPGA_Power_SUSPEND R
  XR58 FPGA_Power_VFS VCC3V3 R
  XR59 FPGA_Power_VBATT VCC3V3 R
  XC243 GND VCC3V3 C
  XC242 GND VCC3V3 C
  XU3 FPGA_Bank_1_2_SPI_CS_N unnamed unnamed GND FPGA_Bank_1_2_SPI_MOSI_CSI_N_MISO0 FPGA_Bank_1_2_SPI_CLK FPGA_Bank_1_2_SPI_D2_MISO3 VCC3V3 W25Q128FVEIG
  XR16 unnamed FPGA_Bank_1_2_SPI_DO_DIN_MISO1 R
  XR17 unnamed FPGA_Bank_1_2_SPI_D1_MISO2 R
  XR20 VCC3V3 unnamed R
  XR19 VCC3V3 unnamed R
  XR18 VCC3V3 FPGA_Bank_1_2_SPI_CS_N R
  XR21 FPGA_Bank_1_2_SPI_D2_MISO3 VCC3V3 R
  XC36 GND VCC3V3 C
  XJP1 FPGA_Bank_1_2_FPGA_M0_CMP_MISO GND JUMPER
  XJP2 FPGA_Bank_1_2_FPGA_M1 GND JUMPER
  XR60 FPGA_Bank_1_2_SD_DAT2 VCC3V3 R
  XR61 FPGA_Bank_1_2_SD_DAT3 VCC3V3 R
  XR62 FPGA_Bank_1_2_SD_CMD VCC3V3 R
  XR63 FPGA_Bank_1_2_SD_DAT0 VCC3V3 R
  XR64 FPGA_Bank_1_2_SD_DAT1 VCC3V3 R
  XC132 GND VCC3V3 C
  XU17 unnamed GND FPGA_Bank_1_2_100MHz VCC3V3 FXO-HC536R
  XR80 VCC3V3 unnamed R
  XC188 GND VCC3V3 C
  XC189 GND FPGA_Bank_1_2_100MHz C
  XU11 FPGA_Bank_1_2_SD_DAT2 GND GND GND FPGA_Bank_1_2_SD_DAT3 FPGA_Bank_1_2_SD_CMD VCC3V3 FPGA_Bank_1_2_SD_CLK GND FPGA_Bank_1_2_SD_DAT0 FPGA_Bank_1_2_SD_DAT1 GND MICRO_SD
  XP3 GND unnamed GND unnamed GND unnamed VCC3V3 GND unnamed GND unnamed GND unnamed GND CONN_7X2
  XR40 VCC3V3 FPGA_Bank_1_2_FPGA_M0_CMP_MISO R
  XR41 FPGA_Bank_1_2_FPGA_M1 VCC3V3 R
  XR76 unnamed FPGA_Power_TMS R
  XR81 unnamed FPGA_Power_TCK R
  XR82 unnamed SPI_Flash_TDO_FPGA_TDO_JTAG R
  XR83 unnamed SPI_Flash_TDO_USB_TDI_FPGA R
  XU26 unnamed GND SPI_Flash_27MHz VCC3V3 FXO-HC536R
  XR86 VCC3V3 unnamed R
  XC241 GND VCC3V3 C
  XC244 GND SPI_Flash_27MHz C
  XP14 unnamed unnamed unnamed FPGA_Bank_0_3_PCIO1 FPGA_Bank_0_3_PCIO2 unnamed FPGA_Bank_0_3_PCIO3 SPI_Flash_RST unnamed unnamed CONN_5X2
  XR93 VCC3V3 unnamed R
  XR118 unnamed FPGA_Bank_0_3_PCIO0 R
  XR116 GND unnamed R
  XR117 FPGA_Bank_0_3_PCIO3 VCC1V5 R
  XR119 unnamed GND R
  XP28 FPGA_Bank_1_2_SD_DAT1 FPGA_Bank_1_2_SD_DAT0 FPGA_Bank_1_2_SD_CLK FPGA_Bank_1_2_SD_CMD FPGA_Bank_1_2_SD_DAT3 FPGA_Bank_1_2_SD_DAT2 VCC3V3 GND CONN_8
  XU1 VCC1V5 DDR3_DDR0_DQ13 DDR3_DDR0_DQ15 DDR3_DDR0_DQ12 VCC1V5 GND GND VCC1V5 GND DDR3_DDR0_UDQS_N DDR3_DDR0_DQ14 GND VCC1V5 DDR3_DDR0_DQ11 DDR3_DDR0_DQ9 DDR3_DDR0_UDQS_P DDR3_DDR0_DQ10 VCC1V5 GND VCC1V5 DDR3_DDR0_UDM DDR3_DDR0_DQ8 GND VCC1V5 GND GND DDR3_DDR0_DQ0 DDR3_DDR0_LDM GND VCC1V5 VCC1V5 DDR3_DDR0_DQ2 DDR3_DDR0_LDQS_P DDR3_DDR0_DQ1 DDR3_DDR0_DQ3 GND GND DDR3_DDR0_DQ6 DDR3_DDR0_LDQS_N VCC1V5 GND GND VTTREF VCC1V5 DDR3_DDR0_DQ4 DDR3_DDR0_DQ7 DDR3_DDR0_DQ5 VCC1V5 unnamed GND DDR3_DDR0_RAS_N DDR3_DDR0_CK_P GND unnamed DDR3_DDR0_ODT VCC1V5 DDR3_DDR0_CAS_N DDR3_DDR0_CK_N VCC1V5 DDR3_DDR0_CKE unnamed unnamed DDR3_DDR0_WE_N DDR3_DDR0_A10 unnamed unnamed GND DDR3_DDR0_BA0 DDR3_DDR0_BA2 unnamed VTTREF GND VCC1V5 DDR3_DDR0_A3 DDR3_DDR0_A0 DDR3_DDR0_A12 DDR3_DDR0_BA1 VCC1V5 GND DDR3_DDR0_A5 DDR3_DDR0_A2 DDR3_DDR0_A1 DDR3_DDR0_A4 GND VCC1V5 DDR3_DDR0_A7 DDR3_DDR0_A9 DDR3_DDR0_A11 DDR3_DDR0_A6 VCC1V5 GND DDR3_DDR0_RESET_N DDR3_DDR0_A13 DDR3_DDR0_A14 DDR3_DDR0_A8 GND MT41J128M16
  XR1 VTTDDR0 DDR3_DDR0_A13 R
  XR10 VTTDDR0 DDR3_DDR0_BA1 VTTDDR0 DDR3_DDR0_A10 VTTDDR0 DDR3_DDR0_WE_N VTTDDR0 DDR3_DDR0_RAS_N RES_NET4
  XR9 VTTDDR0 DDR3_DDR0_A1 VTTDDR0 DDR3_DDR0_A14 VTTDDR0 DDR3_DDR0_A8 VTTDDR0 DDR3_DDR0_A6 RES_NET4
  XR8 VTTDDR0 DDR3_DDR0_BA2 VTTDDR0 DDR3_DDR0_A2 VTTDDR0 DDR3_DDR0_A9 VTTDDR0 DDR3_DDR0_A0 RES_NET4
  XR3 VTTDDR0 DDR3_DDR0_BA0 VTTDDR0 DDR3_DDR0_A5 VTTDDR0 DDR3_DDR0_A7 VTTDDR0 DDR3_DDR0_A3 RES_NET4
  XR2 VTTDDR0 DDR3_DDR0_A11 VTTDDR0 DDR3_DDR0_A4 VTTDDR0 DDR3_DDR0_A12 VTTDDR0 DDR3_DDR0_CAS_N RES_NET4
  XR11 GND unnamed R
  XR12 unnamed GND R
  XC33 VTTREF GND C
  XR4 DDR3_DDR0_CK_N DDR3_DDR0_CK_P R
  XR7 GND DDR3_DDR0_CKE R
  XR6 GND DDR3_DDR0_ODT R
  XR5 GND DDR3_DDR0_RESET_N R
  XC1 VTTDDR0 GND C
  XC2 VTTDDR0 GND C
  XC3 VTTDDR0 GND C
  XC4 VTTDDR0 GND C
  XC5 VTTDDR0 GND C
  XC6 VTTDDR0 GND C
  XC7 VTTDDR0 GND C
  XC8 VTTDDR0 GND C
  XC9 VTTDDR0 GND C
  XC10 VTTDDR0 GND C
  XC11 VTTDDR0 GND C
  XC12 VTTDDR0 GND C
  XC13 VTTDDR0 GND C
  XC14 VTTDDR0 GND C
  XC15 VTTDDR0 GND C
  XC16 GND VCC1V5 C
  XC17 GND VCC1V5 C
  XC18 GND VCC1V5 C
  XC19 GND VCC1V5 C
  XC20 GND VCC1V5 C
  XC21 GND VCC1V5 C
  XC22 GND VCC1V5 C
  XC23 GND VCC1V5 C
  XC24 GND VCC1V5 C
  XC25 GND VCC1V5 C
  XC26 GND VCC1V5 C
  XC27 GND VCC1V5 C
  XC28 GND VCC1V5 C
  XC29 GND VCC1V5 C
  XC30 GND VCC1V5 C
  XC31 GND VCC1V5 C
  XC32 GND VCC1V5 C
  XC174 VTTDDR0 GND C
  XC176 VTTDDR0 GND C
  XC178 VTTDDR0 GND C
  XC180 VTTDDR0 GND C
  XC182 VTTDDR0 GND C
  XC184 VTTDDR0 GND C
  XC186 VTTDDR0 GND C
  XC187 VTTDDR0 GND C
  XC207 VTTDDR0 GND C
  XC209 VTTDDR0 GND C
  XJ8 unnamed unnamed GND unnamed DisplayPort_DPTXCONFIG1 DisplayPort_DPTXCONFIG2 unnamed GND unnamed FPGA_Bank_1_2_DPTXHPD GND GND unnamed unnamed unnamed GND unnamed unnamed GND unnamed DISPLAY_PORT
  XJ9 unnamed unnamed GND unnamed DisplayPort_DPRXCONFIG1 DisplayPort_DPRXCONFIG2 unnamed GND unnamed FPGA_Bank_1_2_DPRXHPD GND GND unnamed unnamed unnamed GND unnamed unnamed GND unnamed DISPLAY_PORT
  XR25 unnamed GND R
  XF3 VCC4V0 unnamed FUSE
  XR42 DisplayPort_DPTXCONFIG1 GND R
  XR43 DisplayPort_DPTXCONFIG2 GND R
  XR45 DisplayPort_DPRXCONFIG1 GND R
  XR46 DisplayPort_DPRXCONFIG2 GND R
  XR47 FPGA_Bank_1_2_DPRXHPD GND R
  XR44 FPGA_Bank_1_2_DPTXHPD GND R
  XD3 unnamed unnamed DIODE
  XF2 VCC4V0 unnamed FUSE
  XD11 unnamed unnamed DIODE
  XC47 unnamed GND C
  XC49 unnamed GND C
  XC264 DisplayPort_DPRX_LANEN3 unnamed C
  XC265 DisplayPort_DPRX_LANEP3 unnamed C
  XC260 DisplayPort_DPRX_LANEN2 unnamed C
  XC261 DisplayPort_DPRX_LANEP2 unnamed C
  XC266 DisplayPort_DPRX_LANEN1 unnamed C
  XC267 DisplayPort_DPRX_LANEP1 unnamed C
  XC262 DisplayPort_DPRX_LANEN0 unnamed C
  XC263 DisplayPort_DPRX_LANEP0 unnamed C
  XC254 DisplayPort_DPTX_LANEP0 unnamed C
  XC255 DisplayPort_DPTX_LANEN0 unnamed C
  XC104 DisplayPort_DPTX_LANEP1 unnamed C
  XC106 DisplayPort_DPTX_LANEN1 unnamed C
  XC256 DisplayPort_DPTX_LANEP2 unnamed C
  XC257 DisplayPort_DPTX_LANEN2 unnamed C
  XC251 DisplayPort_DPTX_LANEP3 unnamed C
  XC253 DisplayPort_DPTX_LANEN3 unnamed C
  XC50 DisplayPort_DPTXAUXCH_P unnamed C
  XC100 DisplayPort_DPTXAUXCH_N unnamed C
  XC258 DisplayPort_DPRXAUXCH_P unnamed C
  XC259 DisplayPort_DPRXAUXCH_N unnamed C
  XR122 unnamed GND R
  XR123 unnamed unnamed R
  XC238 Ethernet_XTAL1_50MHZ GND C
  XL6 VCC3V3 Ethernet_AVDD3V3 INDUCTOR
  XC235 Ethernet_XTAL2_50MHZ GND C
  XR89 unnamed GND R
  XR92 unnamed VCC3V3 R
  XX2 Ethernet_XTAL2_50MHZ Ethernet_XTAL1_50MHZ CRYSTAL
  XC239 VCC3V3 GND C
  XU23 GND GND unnamed GND Ethernet_MAC_SDA Ethernet_MAC_SCL Ethernet_MAC_WP VCC3V3 24AA02E48
  XU20 unnamed unnamed unnamed unnamed Ethernet_ETH_RXCTL Ethernet_ETH_RXD0 Ethernet_ETH_VCC3V3 Ethernet_ETH_RXD1 Ethernet_ETH_RXD2 Ethernet_ETH_RXD3 Ethernet_ETH_RXCLK unnamed Ethernet_ETH_INT_B Ethernet_ETH_VCC3V3 Ethernet_ETH_TXCLK Ethernet_ETH_TXD0 Ethernet_ETH_TXD1 Ethernet_ETH_TXD2 Ethernet_ETH_TXD3 Ethernet_ETH_TXCTL Ethernet_ETH_VCC1V0 Ethernet_ETH_RESET_B Ethernet_ETH_VCC1V0 Ethernet_ETH_MDC Ethernet_ETH_MDIO unnamed unnamed unnamed unnamed Ethernet_ETH_VCC1V0 Ethernet_ETH_VCC3V3 GND unnamed unnamed Ethernet_ETH_VCC1V0 Ethernet_AVDD3V3 Ethernet_XTAL1_50MHZ Ethernet_XTAL2_50MHZ unnamed unnamed unnamed GND unnamed unnamed Ethernet_AVDD3V3 unnamed unnamed Ethernet_ETH_VCC1V0 GND RTL8211E-VL
  XJ6 GND unnamed GND unnamed Ethernet_LED0 Ethernet_LED1 unnamed unnamed unnamed unnamed unnamed unnamed unnamed unnamed unnamed RJ45(HFJ11-1GO1ERL)
  XR71 unnamed VCC3V3 R
  XR70 unnamed Ethernet_LED0 R
  XR69 unnamed GND R
  XR73 unnamed Ethernet_LED1 R
  XR74 unnamed GND R
  XR75 unnamed VCC3V3 R
  XC210 VCC3V3 GND C
  XC217 VCC3V3 GND C
  XC224 Ethernet_AVDD3V3 GND C
  XC227 Ethernet_AVDD3V3 GND C
  XC230 Ethernet_AVDD3V3 GND C
  XL7 VCC3V3 Ethernet_ETH_VCC3V3 INDUCTOR
  XC211 VCC3V3 GND C
  XC218 VCC3V3 GND C
  XC225 Ethernet_ETH_VCC3V3 GND C
  XC228 Ethernet_ETH_VCC3V3 GND C
  XC231 Ethernet_ETH_VCC3V3 GND C
  XL1 Ethernet_VCC1V0 Ethernet_ETH_VCC1V0 INDUCTOR
  XC212 Ethernet_VCC1V0 GND C
  XC223 Ethernet_ETH_VCC1V0 GND C
  XC232 Ethernet_ETH_VCC1V0 GND C
  XC233 Ethernet_ETH_VCC1V0 GND C
  XC234 Ethernet_ETH_VCC1V0 GND C
  XC220 Ethernet_ETH_VCC3V3 GND C
  XC229 Ethernet_ETH_VCC1V0 GND C
  XC226 Ethernet_ETH_VCC1V0 GND C
  XR67 Ethernet_ETH_VCC3V3 Ethernet_ETH_RXD3 R
  XR66 Ethernet_ETH_VCC3V3 Ethernet_ETH_RXD2 R
  XR65 Ethernet_ETH_VCC3V3 Ethernet_ETH_RXD1 R
  XR49 Ethernet_ETH_VCC3V3 Ethernet_ETH_RXD0 R
  XR48 GND Ethernet_ETH_RXCTL R
  XC216 GND Ethernet_ETH_RXCLK C
  XR50 Ethernet_ETH_VCC3V3 Ethernet_ETH_MDIO R
  XR51 Ethernet_ETH_RESET_B VCC3V3 R
  XC222 Ethernet_ETH_RESET_B GND C
  XU19 unnamed VCC3V3 GND Ethernet_VCC1V0 unnamed GND MCP1825
  XR38 unnamed Ethernet_VCC1V0 R
  XR39 GND unnamed R
  XR22 unnamed VCC3V3 R
  XC203 VCC3V3 GND C
  XC204 Ethernet_VCC1V0 GND C
  XC219 Ethernet_ETH_VCC3V3 GND C
  XC214 Ethernet_ETH_VCC3V3 GND C
  XK1 VCC3V3 unnamed GND CONN_3
  XK2 GND unnamed VCC3V3 CONN_3
  XR151 Ethernet_MAC_WP unnamed R
  XU25 GPIOs_PRSNT VCC3V3 FPGA_Bank_0_3_PCIE_RESET GND FPGA_Bank_0_3_DIFFCLK_XP FPGA_Bank_0_3_DIFFCLK_XN GND FPGA_Bank_0_3_DIFFIO_A1P FPGA_Bank_0_3_DIFFIO_A1N GND FPGA_Bank_0_3_DIFFIO_YP VCC12V0 GND FPGA_Bank_0_3_DIFFIO_A2P FPGA_Bank_0_3_DIFFIO_A2N GND GND FPGA_Bank_0_3_DIFFIO_A3P FPGA_Bank_0_3_DIFFIO_A3N GND GND FPGA_Bank_0_3_DIFFCLK_A0P VCC12V0 FPGA_Bank_0_3_DIFFCLK_A0N GND FPGA_Bank_0_3_DIFFIO_ZP unnamed GND FPGA_Bank_0_3_DIFFIO_A4P FPGA_Bank_0_3_DIFFIO_A4N GND GND FPGA_Bank_0_3_DIFFIO_A5P GND FPGA_Bank_0_3_DIFFIO_A5N GND GND FPGA_Bank_0_3_DIFFIO_A6P FPGA_Bank_0_3_DIFFIO_A6N GND GND FPGA_Bank_0_3_DIFFCLK_A1P FPGA_Bank_0_3_DIFFCLK_A1N GND FPGA_Bank_0_3_DIFFIO_A0P FPGA_Bank_0_3_DIFFIO_A0N FPGA_Bank_0_3_DIFFIO_B0P FPGA_Bank_0_3_DIFFIO_B0N VCC3V3 VCC12V0 VCC3V3 FPGA_Bank_0_3_DIFFIO_XN FPGA_Bank_0_3_DIFFIO_YN GND FPGA_Bank_0_3_DIFFIO_B1P FPGA_Bank_0_3_DIFFIO_B1N GND GPIOs_PRSNT GND FPGA_Bank_0_3_DIFFIO_B2P VCC12V0 FPGA_Bank_0_3_DIFFIO_B2N GND GND FPGA_Bank_0_3_DIFFIO_B3P FPGA_Bank_0_3_DIFFIO_B3N GND GND FPGA_Bank_0_3_DIFFCLK_B0P FPGA_Bank_0_3_DIFFCLK_B0N GND VCC12V0 FPGA_Bank_0_3_DIFFIO_ZN GPIOs_PRSNT GND FPGA_Bank_0_3_DIFFIO_B4P FPGA_Bank_0_3_DIFFIO_B4N GND GND FPGA_Bank_0_3_DIFFIO_B5P FPGA_Bank_0_3_DIFFIO_B5N GND GND GND FPGA_Bank_0_3_DIFFIO_B6P FPGA_Bank_0_3_DIFFIO_B6N GND GND FPGA_Bank_0_3_DIFFCLK_B1P FPGA_Bank_0_3_DIFFCLK_B1N GND GPIOs_PRSNT GND FPGA_Bank_0_3_SMCLK FPGA_Bank_0_3_SMDATA GND VCC3V3 FPGA_Bank_0_3_DIFFIO_XP TIMVIDEOS-PCIE-8X
  XC39 VCC3V3 GND C
  XC40 VCC3V3 GND C
  XC41 VCC3V3 GND C
  XC42 VCC3V3 GND C
  XC43 VCC3V3 GND C
  XC44 VCC3V3 GND C
  XC52 VCC3V3 GND C
  XC53 VCC3V3 GND C
  XC62 GND USB_XTALIN C
  XC64 USB_XTALIOUT GND C
  XX1 USB_XTALIOUT USB_XTALIN CRYSTAL
  XR35 unnamed VCC3V3 R
  XR33 USB_U1_SDA VCC3V3 R
  XR34 Ethernet_MAC_SCL VCC3V3 R
  XR36 GND unnamed R
  XU18 VCC3V3 FPGA_Bank_1_2_USB_D6 GND unnamed FPGA_Bank_1_2_USB_D7 GND unnamed unnamed USB_CPEN USB_USB_DP USB_USB_DM FPGA_Bank_1_2_USB_NXT unnamed VCC3V3 unnamed USB_ID unnamed unnamed FPGA_Bank_1_2_USB_REFCLK FPGA_Bank_1_2_USB_RESETB unnamed FPGA_Bank_1_2_USB_STP FPGA_Bank_1_2_USB_D0 unnamed FPGA_Bank_1_2_USB_DIR VCC3V3 GND FPGA_Bank_1_2_USB_D1 FPGA_Bank_1_2_USB_D2 FPGA_Bank_1_2_USB_D3 FPGA_Bank_1_2_USB_D4 GND FPGA_Bank_1_2_USB_D5 USB3340
  XJ1 USB_USB_5V USB_USB_DM USB_USB_DP USB_ID GND USB_MICRO_B
  XU2 VCC3V3 USB_XTALIOUT unnamed USB_XTALIN GND unnamed unnamed unnamed VCC3V3 USB_CYDP USB_CYDN GND GND VCC3V3 GND unnamed FPGA_Bank_1_2_CY_T0 unnamed unnamed FPGA_Bank_1_2_CY_IFCLK unnamed unnamed Ethernet_MAC_SCL FPGA_Bank_1_2_CY_RD0 USB_U1_SDA FPGA_Bank_1_2_CY_RD FPGA_Bank_1_2_CY_WR VCC3V3 FPGA_Bank_1_2_CY_FD0 FPGA_Bank_1_2_CY_FD1 FPGA_Bank_1_2_CY_FD2 FPGA_Bank_1_2_CY_FD3 VCC3V3 GND FPGA_Bank_1_2_CY_RD1 FPGA_Bank_1_2_CY_TXD0 FPGA_Bank_1_2_CY_RXD0 FPGA_Bank_1_2_CY_TXD1 FPGA_Bank_1_2_CY_RXD1 FPGA_Bank_1_2_CY_FD4 FPGA_Bank_1_2_CY_FD5 FPGA_Bank_1_2_CY_FD6 FPGA_Bank_1_2_CY_FD7 GND VCC3V3 FPGA_Bank_1_2_CY_RD2 GND FPGA_Bank_1_2_CY_CTL3 FPGA_Bank_1_2_CY_CTL4 VCC3V3 FPGA_Bank_1_2_CY_CTL0 FPGA_Bank_1_2_CY_CTL1 FPGA_Bank_1_2_CY_CTL2 FPGA_Bank_1_2_CY_PC0 FPGA_Bank_1_2_CY_PC1 FPGA_Bank_1_2_CY_PC2 FPGA_Bank_1_2_CY_RD3 FPGA_Bank_1_2_CY_PC3 FPGA_Bank_1_2_CY_PC4 FPGA_Bank_1_2_CY_PC5 FPGA_Bank_1_2_CY_PC6 FPGA_Bank_1_2_CY_PC7 GND VCC3V3 FPGA_Bank_1_2_CY_PA0 FPGA_Bank_1_2_CY_PA1 FPGA_Bank_1_2_CY_PA2 FPGA_Bank_1_2_CY_RD4 FPGA_Bank_1_2_CY_PA3 FPGA_Bank_1_2_CY_PA4 FPGA_Bank_1_2_CY_PA5 FPGA_Bank_1_2_CY_PA6 FPGA_Bank_1_2_CY_PA7 GND FPGA_Bank_1_2_CY_CTL5 USB_CYP_RESET VCC3V3 unnamed FPGA_Bank_1_2_CY_RD5 FPGA_Bank_1_2_CY_FD8 FPGA_Bank_1_2_CY_FD9 FPGA_Bank_1_2_CY_FD10 FPGA_Bank_1_2_CY_FD11 FPGA_Bank_1_2_CY_INT5 VCC3V3 unnamed unnamed unnamed unnamed VCC3V3 unnamed unnamed unnamed unnamed GND FPGA_Bank_1_2_CY_FD12 FPGA_Bank_1_2_CY_FD13 FPGA_Bank_1_2_CY_FD14 FPGA_Bank_1_2_CY_FD15 GND CY7C68013A_100AC
  XC54 VCC3V3 GND C
  XC58 VCC3V3 GND C
  XC66 VCC3V3 GND C
  XC201 VCC3V3 GND C
  XC202 VCC3V3 GND C
  XR13 GND unnamed R
  XC35 unnamed GND C
  XC34 unnamed GND C
  XR30 unnamed USB_USB_5V R
  XC37 GND unnamed C
  XR14 unnamed SPI_Flash_TDO_FPGA_TDO_JTAG R
  XR23 unnamed SPI_Flash_TDO_USB_TDI_FPGA R
  XR24 unnamed FPGA_Power_TMS R
  XR26 unnamed FPGA_Power_TCK R
  XR15 unnamed FPGA_Power_PROG_B R
  XR28 unnamed FPGA_Power_DONE R
  XR27 unnamed FPGA_Bank_1_2_INIT_B R
  XD2 unnamed GND LED
  XR31 unnamed unnamed R
  XP11 unnamed CONN_1
  XP12 unnamed CONN_1
  XR32 unnamed GND R
  XP13 unnamed CONN_1
  XGS2 unnamed VCC3V3 GS2
  XR37 unnamed GND R
  XU24 USB_USB_5V USB_USB_5V GND unnamed USB_CPEN unnamed unnamed VCC12V0 GND BDXXGA5WEFJ_
  XC240 USB_USB_5V GND C
  XC38 VCC12V0 GND C
  XP17 unnamed USB_CYDN USB_CYDP GND unnamed CONN_5
  XP16 USB_USB_5V USB_USB_DM USB_USB_DP GND unnamed CONN_5
  XP18 USB_U1_SDA Ethernet_MAC_SDA CONN_2
  XR72 USB_CYP_RESET VCC3V3 R
  XC46 USB_CYP_RESET GND C
  XD12 USB_CYP_RESET SPI_Flash_RST DIODESCH
  XD13 FPGA_Power_PROG_B SPI_Flash_RST DIODESCH
  XJ7 unnamed USB_CYDN USB_CYDP GND GND GND USB
  XK3 unnamed FPGA_Bank_1_2_CYPRESS_RESET USB_CYP_RESET CONN_3
  XC191 VCC1V2 GND C
  XC193 VCC1V2 GND C
  XC194 VCC1V2 GND C
  XC195 VCC1V2 GND C
  XC196 VCC1V2 GND C
  XC197 VCC1V2 GND C
  XC198 VCC1V2 GND C
  XC199 VCC1V2 GND C
  XC200 VCC1V2 GND C
  XR85 GND unnamed R
  XC113 VTTREF GND C
  XC192 VTTREF GND C
  XR68 VCC1V2 unnamed R
  XC245 FPGA_Bank_0_3_MGTREFCLK0_101_P unnamed C
  XC246 FPGA_Bank_0_3_MGTREFCLK0_101_N unnamed C
  XC248 FPGA_Bank_0_3_MGT135MHz_P unnamed C
  XC247 FPGA_Bank_0_3_MGT135MHz_N unnamed C
  XU28 GND GND GND unnamed SMA_CON
  XU29 GND GND GND unnamed SMA_CON
  XC250 FPGA_Bank_0_3_MGTSMACLK_N unnamed C
  XC249 FPGA_Bank_0_3_MGTSMACLK_P unnamed C
  XU27 unnamed unnamed GND unnamed unnamed VCC3V3 FXO-LC73
  XR120 unnamed VCC3V3 R
  XP15 VCC3V3 VCC1V5 FPGA_Bank_0_3_DEBUG_IO0 FPGA_Bank_0_3_DEBUG_IO1 GND CONN_5
  XSW1 unnamed GND SW_PUSH
  XR54 FPGA_Bank_0_3_SWITCH unnamed R
  XJ4 FPGA_Bank_1_2_TMDS_RX1_2_P FPGA_Bank_1_2_TMDS_RX1_CLK_P GND FPGA_Bank_1_2_TMDS_RX1_CLK_N HDMI_P1_CEC unnamed HDMI_P1_SCL HDMI_P1_SDA GND unnamed HDMI_P1_HOT GND FPGA_Bank_1_2_TMDS_RX1_2_N FPGA_Bank_1_2_TMDS_RX1_1_P GND FPGA_Bank_1_2_TMDS_RX1_1_N FPGA_Bank_1_2_TMDS_RX1_0_P GND FPGA_Bank_1_2_TMDS_RX1_0_N HDMI
  XU15 HDMI_HDMI_VCC5V0 FPGA_Bank_1_2_TMDS_RX1_0_P GND FPGA_Bank_1_2_TMDS_RX1_0_N FPGA_Bank_1_2_TMDS_RX1_CLK_P GND FPGA_Bank_1_2_TMDS_RX1_CLK_N FPGA_Bank_1_2_TMDS_RX1_CEC FPGA_Bank_1_2_TMDS_RX1_SCL FPGA_Bank_1_2_TMDS_RX1_SDA FPGA_Bank_1_2_TMDS_RX1_HOT VCC3V3 HDMI_P1_HOT HDMI_P1_SDA HDMI_P1_SCL HDMI_P1_CEC FPGA_Bank_1_2_TMDS_RX1_CLK_N GND FPGA_Bank_1_2_TMDS_RX1_CLK_P FPGA_Bank_1_2_TMDS_RX1_0_N GND FPGA_Bank_1_2_TMDS_RX1_0_P GND FPGA_Bank_1_2_TMDS_RX1_1_N GND FPGA_Bank_1_2_TMDS_RX1_1_P FPGA_Bank_1_2_TMDS_RX1_2_N GND FPGA_Bank_1_2_TMDS_RX1_2_P GND unnamed unnamed FPGA_Bank_1_2_TMDS_RX1_2_P GND FPGA_Bank_1_2_TMDS_RX1_2_N FPGA_Bank_1_2_TMDS_RX1_1_P GND FPGA_Bank_1_2_TMDS_RX1_1_N IP4776CZ38
  XC171 unnamed GND C
  XJ3 FPGA_Bank_1_2_TMDS_TX1_2_P FPGA_Bank_1_2_TMDS_TX1_CLK_P GND FPGA_Bank_1_2_TMDS_TX1_CLK_N HDMI_P2_CEC unnamed HDMI_P2_SCL HDMI_P2_SDA GND HDMI_HDMI_TX1_VCC5V0 HDMI_P2_HOT GND FPGA_Bank_1_2_TMDS_TX1_2_N FPGA_Bank_1_2_TMDS_TX1_1_P GND FPGA_Bank_1_2_TMDS_TX1_1_N FPGA_Bank_1_2_TMDS_TX1_0_P GND FPGA_Bank_1_2_TMDS_TX1_0_N HDMI
  XU13 HDMI_HDMI_VCC5V0 FPGA_Bank_1_2_TMDS_TX1_0_P GND FPGA_Bank_1_2_TMDS_TX1_0_N FPGA_Bank_1_2_TMDS_TX1_CLK_P GND FPGA_Bank_1_2_TMDS_TX1_CLK_N FPGA_Bank_1_2_TMDS_TX1_CEC FPGA_Bank_1_2_TMDS_TX1_SCL FPGA_Bank_1_2_TMDS_TX1_SDA FPGA_Bank_1_2_TMDS_TX1_HOT VCC3V3 HDMI_P2_HOT HDMI_P2_SDA HDMI_P2_SCL HDMI_P2_CEC FPGA_Bank_1_2_TMDS_TX1_CLK_N GND FPGA_Bank_1_2_TMDS_TX1_CLK_P FPGA_Bank_1_2_TMDS_TX1_0_N GND FPGA_Bank_1_2_TMDS_TX1_0_P GND FPGA_Bank_1_2_TMDS_TX1_1_N GND FPGA_Bank_1_2_TMDS_TX1_1_P FPGA_Bank_1_2_TMDS_TX1_2_N GND FPGA_Bank_1_2_TMDS_TX1_2_P GND unnamed unnamed FPGA_Bank_1_2_TMDS_TX1_2_P GND FPGA_Bank_1_2_TMDS_TX1_2_N FPGA_Bank_1_2_TMDS_TX1_1_P GND FPGA_Bank_1_2_TMDS_TX1_1_N IP4776CZ38
  XC169 unnamed GND C
  XJ2 FPGA_Bank_1_2_TMDS_TX2_2_P FPGA_Bank_1_2_TMDS_TX2_CLK_P GND FPGA_Bank_1_2_TMDS_TX2_CLK_N HDMI_P4_CEC unnamed HDMI_P4_SCL HDMI_P4_SDA GND HDMI_HDMI_TX2_VCC5V0 HDMI_P4_HOT GND FPGA_Bank_1_2_TMDS_TX2_2_N FPGA_Bank_1_2_TMDS_TX2_1_P GND FPGA_Bank_1_2_TMDS_TX2_1_N FPGA_Bank_1_2_TMDS_TX2_0_P GND FPGA_Bank_1_2_TMDS_TX2_0_N HDMI
  XC170 unnamed GND C
  XR138 HDMI_HDMI_VCC5V0 HDMI_P4_SDA R
  XR140 HDMI_HDMI_VCC5V0 HDMI_P4_SCL R
  XR129 VCC3V3 FPGA_Bank_1_2_TMDS_TX2_SCL R
  XR133 VCC3V3 FPGA_Bank_1_2_TMDS_TX2_SDA R
  XJ5 FPGA_Bank_1_2_TMDS_RX2_2_P FPGA_Bank_1_2_TMDS_RX2_CLK_P GND FPGA_Bank_1_2_TMDS_RX2_CLK_N HDMI_P3_CEC unnamed HDMI_P3_SCL HDMI_P3_SDA GND unnamed HDMI_P3_HOT GND FPGA_Bank_1_2_TMDS_RX2_2_N FPGA_Bank_1_2_TMDS_RX2_1_P GND FPGA_Bank_1_2_TMDS_RX2_1_N FPGA_Bank_1_2_TMDS_RX2_0_P GND FPGA_Bank_1_2_TMDS_RX2_0_N HDMI
  XU21 HDMI_HDMI_VCC5V0 FPGA_Bank_1_2_TMDS_RX2_0_P GND FPGA_Bank_1_2_TMDS_RX2_0_N FPGA_Bank_1_2_TMDS_RX2_CLK_P GND FPGA_Bank_1_2_TMDS_RX2_CLK_N FPGA_Bank_1_2_TMDS_RX2_CEC FPGA_Bank_1_2_TMDS_RX2_SCL FPGA_Bank_1_2_TMDS_RX2_SDA FPGA_Bank_1_2_TMDS_RX2_HOT VCC3V3 HDMI_P3_HOT HDMI_P3_SDA HDMI_P3_SCL HDMI_P3_CEC FPGA_Bank_1_2_TMDS_RX2_CLK_N GND FPGA_Bank_1_2_TMDS_RX2_CLK_P FPGA_Bank_1_2_TMDS_RX2_0_N GND FPGA_Bank_1_2_TMDS_RX2_0_P GND FPGA_Bank_1_2_TMDS_RX2_1_N GND FPGA_Bank_1_2_TMDS_RX2_1_P FPGA_Bank_1_2_TMDS_RX2_2_N GND FPGA_Bank_1_2_TMDS_RX2_2_P GND unnamed unnamed FPGA_Bank_1_2_TMDS_RX2_2_P GND FPGA_Bank_1_2_TMDS_RX2_2_N FPGA_Bank_1_2_TMDS_RX2_1_P GND FPGA_Bank_1_2_TMDS_RX2_1_N IP4776CZ38
  XC179 unnamed GND C
  XR126 VCC3V3 FPGA_Bank_1_2_TMDS_TX2_CEC R
  XR149 GND HDMI_P4_HOT R
  XR144 VCC3V3 HDMI_P4_CEC R
  XR130 VCC3V3 FPGA_Bank_1_2_TMDS_TX1_SDA R
  XR134 VCC3V3 FPGA_Bank_1_2_TMDS_TX1_SCL R
  XR127 VCC3V3 FPGA_Bank_1_2_TMDS_TX1_CEC R
  XR137 HDMI_HDMI_VCC5V0 HDMI_P2_SDA R
  XR139 HDMI_HDMI_VCC5V0 HDMI_P2_SCL R
  XR148 GND HDMI_P2_HOT R
  XR143 VCC3V3 HDMI_P2_CEC R
  XR135 VCC3V3 FPGA_Bank_1_2_TMDS_RX1_SCL R
  XR136 VCC3V3 FPGA_Bank_1_2_TMDS_RX1_SDA R
  XR132 VCC3V3 FPGA_Bank_1_2_TMDS_RX1_CEC R
  XR141 HDMI_HDMI_VCC5V0 HDMI_P1_SDA R
  XR142 HDMI_HDMI_VCC5V0 HDMI_P1_SCL R
  XR146 VCC3V3 HDMI_P1_CEC R
  XR196 HDMI_HDMI_VCC5V0 HDMI_P3_SDA R
  XR197 HDMI_HDMI_VCC5V0 HDMI_P3_SCL R
  XR199 VCC3V3 HDMI_P3_CEC R
  XR193 VCC3V3 FPGA_Bank_1_2_TMDS_RX2_SCL R
  XR194 VCC3V3 FPGA_Bank_1_2_TMDS_RX2_SDA R
  XR192 VCC3V3 FPGA_Bank_1_2_TMDS_RX2_CEC R
  XR125 FPGA_Bank_1_2_TMDS_RX1_0_P VCC3V3 R
  XR128 FPGA_Bank_1_2_TMDS_RX1_1_P VCC3V3 R
  XR131 FPGA_Bank_1_2_TMDS_RX1_2_P VCC3V3 R
  XR124 FPGA_Bank_1_2_TMDS_RX1_CLK_P VCC3V3 R
  XR147 FPGA_Bank_1_2_TMDS_RX1_0_N VCC3V3 R
  XR150 FPGA_Bank_1_2_TMDS_RX1_1_N VCC3V3 R
  XR152 FPGA_Bank_1_2_TMDS_RX1_2_N VCC3V3 R
  XR145 FPGA_Bank_1_2_TMDS_RX1_CLK_N VCC3V3 R
  XR189 FPGA_Bank_1_2_TMDS_RX2_1_P VCC3V3 R
  XR190 FPGA_Bank_1_2_TMDS_RX2_0_P VCC3V3 R
  XR191 FPGA_Bank_1_2_TMDS_RX2_CLK_P VCC3V3 R
  XR188 FPGA_Bank_1_2_TMDS_RX2_2_P VCC3V3 R
  XR201 VCC3V3 FPGA_Bank_1_2_TMDS_RX2_0_N R
  XR200 VCC3V3 FPGA_Bank_1_2_TMDS_RX2_1_N R
  XR198 VCC3V3 FPGA_Bank_1_2_TMDS_RX2_2_N R
  XR203 VCC3V3 FPGA_Bank_1_2_TMDS_RX2_CLK_N R
  XU14 HDMI_HDMI_VCC5V0 FPGA_Bank_1_2_TMDS_TX2_0_P GND FPGA_Bank_1_2_TMDS_TX2_0_N FPGA_Bank_1_2_TMDS_TX2_CLK_P GND FPGA_Bank_1_2_TMDS_TX2_CLK_N FPGA_Bank_1_2_TMDS_TX2_CEC FPGA_Bank_1_2_TMDS_TX2_SCL FPGA_Bank_1_2_TMDS_TX2_SDA FPGA_Bank_1_2_TMDS_TX2_HOT VCC3V3 HDMI_P4_HOT HDMI_P4_SDA HDMI_P4_SCL HDMI_P4_CEC FPGA_Bank_1_2_TMDS_TX2_CLK_N GND FPGA_Bank_1_2_TMDS_TX2_CLK_P FPGA_Bank_1_2_TMDS_TX2_0_N GND FPGA_Bank_1_2_TMDS_TX2_0_P GND FPGA_Bank_1_2_TMDS_TX2_1_N GND FPGA_Bank_1_2_TMDS_TX2_1_P FPGA_Bank_1_2_TMDS_TX2_2_N GND FPGA_Bank_1_2_TMDS_TX2_2_P GND unnamed unnamed FPGA_Bank_1_2_TMDS_TX2_2_P GND FPGA_Bank_1_2_TMDS_TX2_2_N FPGA_Bank_1_2_TMDS_TX2_1_P GND FPGA_Bank_1_2_TMDS_TX2_1_N IP4776CZ38
  XC172 GND HDMI_P1_HOT C
  XR153 HDMI_HDMI_VCC5V0 HDMI_P1_HOT R
  XR205 HDMI_HDMI_VCC5V0 HDMI_P3_HOT R
  XC185 GND HDMI_P3_HOT C
  XU16 HDMI_HDMI_TX1_VCC5V0 GND VCC12V0 ΜA78L00
  XC173 VCC12V0 GND C
  XC175 HDMI_HDMI_TX1_VCC5V0 GND C
  XR195 HDMI_HDMI_TX1_VCC5V0 GND R
  XU22 HDMI_HDMI_TX2_VCC5V0 GND VCC12V0 ΜA78L00
  XC177 VCC12V0 GND C
  XC181 HDMI_HDMI_TX2_VCC5V0 GND C
  XR202 HDMI_HDMI_TX2_VCC5V0 GND R
  XR84 GND unnamed R
  XR88 GND unnamed R
  XP7 FPGA_Bank_1_2_TMDS_RX1_SDA CONN_1
  XP8 FPGA_Bank_1_2_TMDS_RX1_SCL CONN_1
  XP9 FPGA_Bank_1_2_TMDS_RX2_SDA CONN_1
  XP10 FPGA_Bank_1_2_TMDS_RX2_SCL CONN_1
  XP5 FPGA_Bank_1_2_TMDS_TX1_SDA CONN_1
  XP6 FPGA_Bank_1_2_TMDS_TX1_SCL CONN_1
  XP2 FPGA_Bank_1_2_TMDS_TX2_SDA CONN_1
  XP4 FPGA_Bank_1_2_TMDS_TX2_SCL CONN_1
  XC205 HDMI_HDMI_TX1_VCC5V0 GND C
  XC252 HDMI_HDMI_TX2_VCC5V0 GND C
  XU30 HDMI_HDMI_VCC5V0 GND VCC12V0 ΜA78L00
  XC183 VCC12V0 GND C
  XC208 HDMI_HDMI_VCC5V0 GND C
  XR121 HDMI_HDMI_VCC5V0 GND R
  XC206 HDMI_HDMI_VCC5V0 GND C
  XP24 FPGA_Bank_1_2_TMDS_RX1_HOT CONN_1
  XP19 FPGA_Bank_1_2_TMDS_RX1_CEC CONN_1
  XP25 FPGA_Bank_1_2_TMDS_RX2_CEC CONN_1
  XP26 FPGA_Bank_1_2_TMDS_RX2_HOT CONN_1
  XP20 FPGA_Bank_1_2_TMDS_TX1_CEC CONN_1
  XP21 FPGA_Bank_1_2_TMDS_TX1_HOT CONN_1
  XP23 FPGA_Bank_1_2_TMDS_TX2_HOT CONN_1
  XP22 FPGA_Bank_1_2_TMDS_TX2_CEC CONN_1
.ends HDMI2USB

*--- Subcircuit Definitions ---
.subckt TPS54625 1 10 11 12 13 14 15 2 3 4 5 6 7 8 9
* Stub for TPS54625
.ends

.subckt C 1 2
* Stub for C
.ends

.subckt INDUCTOR 1 2
* Stub for INDUCTOR
.ends

.subckt R 1 2
* Stub for R
.ends

.subckt TPS53319 1 10 11 12 13 14 15 16 17 18 19 2 20 21 22 23 3 4 5 6 7 8 9
* Stub for TPS53319
.ends

.subckt CONN_2 1 2
* Stub for CONN_2
.ends

.subckt TPS54560 1 2 3 4 5 6 7 8 9
* Stub for TPS54560
.ends

.subckt GBU15005-G 1 2 3 4
* Stub for GBU15005-G
.ends

.subckt DIODE 1 2
* Stub for DIODE
.ends

.subckt BARREL_JACK 1 2 3
* Stub for BARREL_JACK
.ends

.subckt DIODESCH 1 2
* Stub for DIODESCH
.ends

.subckt FUSE 1 2
* Stub for FUSE
.ends

.subckt TPS51200 1 10 11 2 3 4 5 6 7 8 9
* Stub for TPS51200
.ends

.subckt LED 1 2
* Stub for LED
.ends

.subckt ATX_POWER_SUPPLY 1 2 3 4 5 6
* Stub for ATX_POWER_SUPPLY
.ends

.subckt XC6SLX150T A1 A10 A11 A12 A13 A14 A15 A16 A17 A18 A19 A2 A20 A21 A22 A3 A4 A5 A6 A7 A8 A9 AA1 AA10 AA11 AA12 AA13 AA14 AA15 AA16 AA17 AA18 AA19 AA2 AA20 AA21 AA22 AA3 AA4 AA5 AA6 AA7 AA8 AA9 AB1 AB10 AB11 AB12 AB13 AB14 AB15 AB16 AB17 AB18 AB19 AB2 AB20 AB21 AB22 AB3 AB4 AB5 AB6 AB7 AB8 AB9 B1 B10 B11 B12 B13 B14 B15 B16 B17 B18 B19 B2 B20 B21 B22 B3 B4 B5 B6 B7 B8 B9 C1 C10 C11 C12 C13 C14 C15 C16 C17 C18 C19 C2 C20 C21 C22 C3 C4 C5 C6 C7 C8 C9 D1 D10 D11 D12 D13 D14 D15 D16 D17 D18 D19 D2 D20 D21 D22 D3 D4 D5 D6 D7 D8 D9 E1 E10 E11 E12 E13 E14 E15 E16 E17 E18 E19 E2 E20 E21 E22 E3 E4 E5 E6 E7 E8 E9 F1 F10 F11 F12 F13 F14 F15 F16 F17 F18 F19 F2 F20 F21 F22 F3 F4 F5 F6 F7 F8 F9 G1 G10 G11 G12 G13 G14 G15 G16 G17 G18 G19 G2 G20 G21 G22 G3 G4 G5 G6 G7 G8 G9 H1 H10 H11 H12 H13 H14 H15 H16 H17 H18 H19 H2 H20 H21 H22 H3 H4 H5 H6 H7 H8 H9 J1 J10 J11 J12 J13 J14 J15 J16 J17 J18 J19 J2 J20 J21 J22 J3 J4 J5 J6 J7 J8 J9 K1 K10 K11 K12 K13 K14 K15 K16 K17 K18 K19 K2 K20 K21 K22 K3 K4 K5 K6 K7 K8 K9 L1 L10 L11 L12 L13 L14 L15 L16 L17 L18 L19 L2 L20 L21 L22 L3 L4 L5 L6 L7 L8 L9 M1 M10 M11 M12 M13 M14 M15 M16 M17 M18 M19 M2 M20 M21 M22 M3 M4 M5 M6 M7 M8 M9 N1 N10 N11 N12 N13 N14 N15 N16 N17 N18 N19 N2 N20 N21 N22 N3 N4 N5 N6 N7 N8 N9 P1 P10 P11 P12 P13 P14 P15 P16 P17 P18 P19 P2 P20 P21 P22 P3 P4 P5 P6 P7 P8 P9 R1 R10 R11 R12 R13 R14 R15 R16 R17 R18 R19 R2 R20 R21 R22 R3 R4 R5 R6 R7 R8 R9 T1 T10 T11 T12 T13 T14 T15 T16 T17 T18 T19 T2 T20 T21 T22 T3 T4 T5 T6 T7 T8 T9 U1 U10 U11 U12 U13 U14 U15 U16 U17 U18 U19 U2 U20 U21 U22 U3 U4 U5 U6 U7 U8 U9 V1 V10 V11 V12 V13 V14 V15 V16 V17 V18 V19 V2 V20 V21 V22 V3 V4 V5 V6 V7 V8 V9 W1 W10 W11 W12 W13 W14 W15 W16 W17 W18 W19 W2 W20 W21 W22 W3 W4 W5 W6 W7 W8 W9 Y1 Y10 Y11 Y12 Y13 Y14 Y15 Y16 Y17 Y18 Y19 Y2 Y20 Y21 Y22 Y3 Y4 Y5 Y6 Y7 Y8 Y9
* Stub for XC6SLX150T
.ends

.subckt W25Q128FVEIG 1 2 3 4 5 6 7 8
* Stub for W25Q128FVEIG
.ends

.subckt JUMPER 1 2
* Stub for JUMPER
.ends

.subckt FXO-HC536R 1 2 3 4
* Stub for FXO-HC536R
.ends

.subckt MICRO_SD 1 10 11 12 2 3 4 5 6 7 8 9
* Stub for MICRO_SD
.ends

.subckt CONN_7X2 1 10 11 12 13 14 2 3 4 5 6 7 8 9
* Stub for CONN_7X2
.ends

.subckt CONN_5X2 1 10 2 3 4 5 6 7 8 9
* Stub for CONN_5X2
.ends

.subckt CONN_8 1 2 3 4 5 6 7 8
* Stub for CONN_8
.ends

.subckt MT41J128M16 A1 A2 A3 A7 A8 A9 B1 B2 B3 B7 B8 B9 C1 C2 C3 C7 C8 C9 D1 D2 D3 D7 D8 D9 E1 E2 E3 E7 E8 E9 F1 F2 F3 F7 F8 F9 G1 G2 G3 G7 G8 G9 H1 H2 H3 H7 H8 H9 J1 J2 J3 J7 J8 J9 K1 K2 K3 K7 K8 K9 L1 L2 L3 L7 L8 L9 M1 M2 M3 M7 M8 M9 N1 N2 N3 N7 N8 N9 P1 P2 P3 P7 P8 P9 R1 R2 R3 R7 R8 R9 T1 T2 T3 T7 T8 T9
* Stub for MT41J128M16
.ends

.subckt RES_NET4 1 2 3 4 5 6 7 8
* Stub for RES_NET4
.ends

.subckt DISPLAY_PORT 1 10 11 12 13 14 15 16 17 18 19 2 20 3 4 5 6 7 8 9
* Stub for DISPLAY_PORT
.ends

.subckt CRYSTAL 1 2
* Stub for CRYSTAL
.ends

.subckt 24AA02E48 1 2 3 4 5 6 7 8
* Stub for 24AA02E48
.ends

.subckt RTL8211E-VL 1 10 11 12 13 14 15 16 17 18 19 2 20 21 22 23 24 25 26 27 28 29 3 30 31 32 33 34 35 36 37 38 39 4 40 41 42 43 44 45 46 47 48 5 6 7 8 9 P
* Stub for RTL8211E-VL
.ends

.subckt RJ45(HFJ11-1GO1ERL) 0 1 10 11 12 13 14 2 3 4 5 6 7 8 9
* Stub for RJ45(HFJ11-1GO1ERL)
.ends

.subckt MCP1825 1 2 3 4 5 6
* Stub for MCP1825
.ends

.subckt CONN_3 1 2 3
* Stub for CONN_3
.ends

.subckt TIMVIDEOS-PCIE-8X A1 A10 A11 A12 A13 A14 A15 A16 A17 A18 A19 A2 A20 A21 A22 A23 A24 A25 A26 A27 A28 A29 A3 A30 A31 A32 A33 A34 A35 A36 A37 A38 A39 A4 A40 A41 A42 A43 A44 A45 A46 A47 A48 A49 A5 A6 A7 A8 A9 B1 B10 B11 B12 B13 B14 B15 B16 B17 B18 B19 B2 B20 B21 B22 B23 B24 B25 B26 B27 B28 B29 B3 B30 B31 B32 B33 B34 B35 B36 B37 B38 B39 B4 B40 B41 B42 B43 B44 B45 B46 B47 B48 B49 B5 B6 B7 B8 B9
* Stub for TIMVIDEOS-PCIE-8X
.ends

.subckt USB3340 1 10 11 12 13 14 15 16 17 18 19 2 20 21 22 23 24 25 26 27 28 29 3 30 31 32 33 4 5 6 7 8 9
* Stub for USB3340
.ends

.subckt USB_MICRO_B 1 2 3 4 5
* Stub for USB_MICRO_B
.ends

.subckt CY7C68013A_100AC 1 10 100 11 12 13 14 15 16 17 18 19 2 20 21 22 23 24 25 26 27 28 29 3 30 31 32 33 34 35 36 37 38 39 4 40 41 42 43 44 45 46 47 48 49 5 50 51 52 53 54 55 56 57 58 59 6 60 61 62 63 64 65 66 67 68 69 7 70 71 72 73 74 75 76 77 78 79 8 80 81 82 83 84 85 86 87 88 89 9 90 91 92 93 94 95 96 97 98 99
* Stub for CY7C68013A_100AC
.ends

.subckt CONN_1 1
* Stub for CONN_1
.ends

.subckt GS2 1 2
* Stub for GS2
.ends

.subckt BDXXGA5WEFJ_ 1 2 3 4 5 6 7 8 9
* Stub for BDXXGA5WEFJ_
.ends

.subckt CONN_5 1 2 3 4 5
* Stub for CONN_5
.ends

.subckt USB 1 2 3 4 5 6
* Stub for USB
.ends

.subckt SMA_CON 1 2
* Stub for SMA_CON
.ends

.subckt FXO-LC73 1 2 3 4 5 6
* Stub for FXO-LC73
.ends

.subckt SW_PUSH 1 2
* Stub for SW_PUSH
.ends

.subckt HDMI 1 10 11 12 13 14 15 16 17 18 19 2 3 4 5 6 7 8 9
* Stub for HDMI
.ends

.subckt IP4776CZ38 1 10 11 12 13 14 15 16 17 18 19 2 20 21 22 23 24 25 26 27 28 29 3 30 31 32 33 34 35 36 37 38 4 5 6 7 8 9
* Stub for IP4776CZ38
.ends

.subckt ΜA78L00 1 2 3
* Stub for ΜA78L00
.ends

