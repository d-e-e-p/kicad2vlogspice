* Spice Netlist (renamed)

*--- Top Level ---
.subckt kicad-pyspice-example 
.ends kicad-pyspice-example

