* Spice Netlist (renamed)

*--- Top Level ---
.subckt div 
.ends div

*--- Subcircuit Definitions ---
