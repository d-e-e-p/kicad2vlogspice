* Spice Netlist (renamed)

*--- Top Level ---
.subckt components 
.ends components

